LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.std_logic_signed.all;
USE IEEE.numeric_std.ALL;

PACKAGE HDC_pkg IS
  TYPE vector_of_std_logic_vector2880 IS ARRAY (NATURAL RANGE <>) OF std_logic_vector(2879 DOWNTO 0);
  TYPE class_vector IS ARRAY (0 TO 2879) OF std_logic_vector(6 DOWNTO 0); --max for each bin would be 80 (because 80 samples) so 7 bits
  TYPE bins_sim IS ARRAY (0 TO 29999) OF std_logic_vector(6 DOWNTO 0);
  TYPE class_sim IS ARRAY (0 TO 79) OF integer range 1 to 4;
END HDC_pkg;

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.std_logic_signed.all;
USE IEEE.numeric_std.ALL;
USE work.HDC_pkg.ALL;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY AudioHDC IS
   PORT ( 
			 SW					: IN 	  STD_LOGIC ;
			 CLOCK_50				: IN    STD_LOGIC;
          		 RESET		                        : IN    STD_LOGIC;
			 START_BIT                       	: OUT   STD_LOGIC; 
			 DONE_BIT				: OUT   STD_LOGIC;
			 PRED_LIGHT                       	: OUT   STD_LOGIC_VECTOR(3 DOWNTO 0);
			 TESTS		                       	: OUT   STD_LOGIC_VECTOR (4 DOWNTO 0);
			 CORRECT_HEXONE				: OUT	  STD_LOGIC_VECTOR (6 DOWNTO 0);
			 CORRECT_HEXTWO				: OUT	  STD_LOGIC_VECTOR (6 DOWNTO 0));
END AudioHDC;


ARCHITECTURE Behavior OF AudioHDC IS
  
  
--  component lpmDiv
--	PORT
--	(
--		clock		: IN STD_LOGIC ;
--		denom		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
--		numer		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
--		quotient	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
--		remain		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
--	);
--  END component;

  
--  component DivFunction
--		PORT(
--		clk    : in  std_logic;             --    clk.clk
--		areset : in  std_logic;             -- areset.reset
--		en     : in  std_logic_vector(0 downto 0); --     en.en
--		a      : in  std_logic_vector(31 downto 0); --      a.a
--		b      : in  std_logic_vector(31 downto 0); --      b.b
--		q      : out std_logic_vector(31 downto 0)                     --      q.q
--	);
--  END component;
	
  component Bins_ROM
		port(
			address				: IN STD_LOGIC_VECTOR (14  DOWNTO 0);
			clock				: IN STD_LOGIC;
			q				: OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
		);
  end component;
  component posHV_RAM
		port(
  		clock					: IN STD_LOGIC;
		data					: IN STD_LOGIC_VECTOR (2879 DOWNTO 0);
		rdaddress				: IN STD_LOGIC_VECTOR (6 DOWNTO 0);
		rden					: IN STD_LOGIC;
		wraddress				: IN STD_LOGIC_VECTOR (6 DOWNTO 0);
		wren					: IN STD_LOGIC;
		q					: OUT STD_LOGIC_VECTOR (2879 DOWNTO 0)
		);
  end component;
  

  component levHV_RAM
		port(
  		clock					: IN STD_LOGIC;
		data					: IN STD_LOGIC_VECTOR (2879 DOWNTO 0);
		rdaddress				: IN STD_LOGIC_VECTOR (6 DOWNTO 0);
		rden					: IN STD_LOGIC;
		wraddress				: IN STD_LOGIC_VECTOR (6 DOWNTO 0);
		wren					: IN STD_LOGIC;
		q					: OUT STD_LOGIC_VECTOR (2879 DOWNTO 0)
		);
  end component;
  
--  component col_sum_RAM 
--		PORT(
--		clock					: IN STD_LOGIC  := '1';
--		data					: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
--		rdaddress				: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
--		wraddress				: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
--		wren					: IN STD_LOGIC  := '0';
--		q					: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
--	);
--	end component col_sum_RAM;
  
  COMPONENT rng_xoshiro128plusplus
     generic (
        -- Default seed value.
        init_seed:  std_logic_vector(127 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
        -- Enable optional pipeline stage in output calculation.
        -- This uses an extra 32-bit register but tends to improve
        -- the timing performance of the circuit.
        -- If the pipeline stage is enabled, two clock cycles are needed
        -- before valid output appears after reset and after re-seeding.
        -- If the pipeline stage is disabled, just one clock cycle is needed.
        pipeline:   boolean := true );
	  PORT(	  
		  -- Clock, rising edge active.
        clk:        in  std_logic;
        -- Synchronous reset, active high.
        rst:        in  std_logic;
        -- High to request re-seeding of the generator.
        reseed:     in  std_logic;
        -- New seed value (must be valid when reseed = '1').
        newseed:    in  std_logic_vector(127 downto 0);
        -- High when the user accepts the current random data word
        -- and requests new random data for the next clock cycle.
        out_ready:  in  std_logic;
        -- High when valid random data is available on the output.
        -- This signal is low for 1 or 2 clock cycles after reset and
        -- after re-seeding, and high in all other cases.
        out_valid:  out std_logic;
        -- Random output data (valid when out_valid = '1').
        -- A new random word appears after every rising clock edge
        -- where out_ready = '1'.
        out_data:   out std_logic_vector(31 downto 0) );
  END COMPONENT;
  
  TYPE state IS (START, POSITION_HVS, HV_SETUP, HV_STORE, HV_READY, LEV_HV_FIRST, LEVEL_HVS, LEVEL_HV_FLIP, LEVEL_HV_SET, TRAIN, AUDIO_ENC, ENC_BIN_SETUP, ENC_BIN_SET, ENC_BIN_VAL, AUDIO_ENC_TEST, TEST_BIN_VEC, INF, INF_RES, RETRAIN, RESULT);
  SIGNAL Mealy_state: state;
  
  --for sim
  --constant binsconst : bins_sim := ("0000000", "0010100", "0000000", "0000000", "0000000", "0000000", "0001010", "0000101", "0001111", "0001010", "0000101", "0001010", "0001111", "0000101", "0001111", "0000101", "0011110", "0001111", "0010100", "0000101", "0010100", "0000101", "0000101", "0000101", "0001111", "0000101", "0000101", "0000101", "0011001", "0000101", "0000101", "0100011", "0011110", "0000000", "0000101", "0000000", "0000000", "0000000", "0000101", "0000000", "0000000", "0000000", "0000000", "0001111", "0000000", "0000000", "0001010", "0101000", "0001111", "0101000", "0000101", "0000101", "0000101", "0001111", "0001010", "0001010", "0000101", "0011001", "0101000", "0100011", "0000101", "0000101", "0000101", "0000101", "0000101", "0000000", "0000101", "0000000", "0000000", "0000101", "0001010", "0010100", "0011001", "0100011", "0101000", "0011001", "0000000", "0000101", "0000101", "0000000", "0011110", "0000101", "0000000", "0100011", "0000101", "0001010", "0000101", "0001010", "0000101", "0000000", "0010100", "0011001", "0101101", "0000000", "0101101", "0100011", "0100011", "0000000", "0000101", "0000101", "0100000", "0110000", "0100001", "0010001", "0001100", "0100011", "0100100", "0100010", "0100000", "0010010", "0100001", "0010111", "0011111", "0101010", "0100100", "0011011", "1000000", "0011010", "0011101", "0011010", "0100000", "0010010", "0001011", "0100001", "0100001", "0101000", "0010110", "0010110", "0101000", "0001110", "0011010", "0100010", "0011110", "0010101", "0111001", "0110011", "0011101", "0101011", "0100100", "0001010", "0001011", "0100101", "0010000", "0111100", "0001011", "0010100", "0011111", "0100110", "0010110", "0100000", "0010000", "0011101", "0010011", "0010110", "0011111", "0010110", "0000111", "0100001", "0100010", "0011000", "0010101", "0101010", "0101110", "0011010", "0100010", "0101001", "0010101", "0011001", "0001001", "0001101", "0101001", "0101011", "0101111", "0110001", "0110011", "0100010", "0011100", "0101000", "0100100", "0001000", "0110111", "0110101", "0010111", "0111000", "0101110", "0010010", "0011000", "0110011", "0011101", "0001101", "0100110", "0011111", "1000101", "0001101", "0110000", "0101100", "0100011", "0011111", "0110101", "0110100", "0101101", "0111110", "0101101", "0011000", "0010000", "0101110", "0101001", "0100101", "0100100", "0010100", "0100110", "0011001", "0101000", "0101100", "0011110", "0011110", "1000100", "0011100", "0100011", "0010000", "0100011", "0010100", "0001100", "0100011", "0100100", "0101010", "0011011", "0010011", "0100011", "0001101", "0011101", "0100111", "0100101", "0001110", "0100101", "0100100", "0100011", "0110100", "0101111", "0001001", "0001010", "0100101", "0010001", "0111110", "0001110", "0011001", "0100011", "0101010", "0011000", "0100011", "0010011", "0100001", "0010110", "0011110", "0100011", "0011010", "0001000", "0100111", "0101110", "0100000", "0011100", "0101001", "0011100", "0001111", "0100001", "0101000", "0010101", "0100010", "0001100", "0001111", "0101010", "0101110", "0110001", "0110011", "0110110", "0100110", "0011101", "0101000", "0100100", "0001010", "0110110", "0110101", "0011000", "0111000", "0111001", "0010001", "0011111", "0110101", "0011101", "0001110", "0100000", "0011000", "0111100", "0010010", "0111001", "0110100", "0101001", "0011010", "0100110", "0100101", "0001101", "0011001", "0001111", "0010000", "0001011", "0100010", "0101001", "0100110", "0100110", "0010100", "0100111", "0011011", "0110011", "0101110", "0100001", "0100001", "0111101", "0011110", "0100011", "0010011", "0100001", "0010011", "0001101", "0100001", "0011000", "0101000", "0100011", "0011001", "0101101", "0010001", "0010111", "0011111", "0100000", "0011001", "1000001", "0111110", "0011011", "0101000", "0100101", "0010000", "0010000", "0111110", "0010100", "0110010", "0010010", "0100010", "0110000", "0111111", "0100011", "0110110", "0011011", "0101101", "0100001", "0100100", "0100110", "0011011", "0001001", "0101111", "0110010", "0100111", "0100001", "0111110", "0100111", "0010110", "0011110", "0100001", "0010001", "0101100", "0001101", "0010101", "0010100", "0010101", "0010110", "0010101", "0011000", "0010001", "0001100", "0010001", "0010000", "0001101", "0011000", "0011101", "0001100", "0010110", "0010110", "0001000", "0100111", "0010010", "0001010", "0000110", "0010011", "0010001", "0100110", "0010110", "0010001", "0010001", "0001110", "0010001", "0011011", "0011011", "0000010", "0001000", "0000011", "0000011", "0000010", "0000110", "0001010", "0001000", "0000111", "0000100", "0001001", "0000101", "0101101", "0001001", "0001000", "0000110", "0010110", "0000101", "0000111", "0010000", "0000110", "0000011", "0000011", "0000110", "0001000", "0001001", "0011110", "0000101", "0001010", "0000100", "0001000", "0001001", "0001001", "0000011", "0000111", "0000111", "0001000", "0001100", "0001100", "0000100", "0000100", "0010001", "0011001", "0100000", "0001111", "0011101", "0100111", "0110100", "0011011", "0101011", "0011000", "0100111", "0011100", "0011111", "0110000", "0011111", "0001100", "0111001", "1000000", "0101111", "0011110", "0111011", "0100011", "0010101", "0110111", "1000010", "0011111", "0110010", "0001110", "0010111", "0000011", "0000100", "0000100", "0000100", "0000100", "0000011", "0000011", "0000011", "0000100", "0001011", "0000100", "0001100", "0000100", "0000101", "0001011", "0000010", "0100001", "0000100", "0000011", "0000011", "0000011", "0000110", "0010101", "0010100", "0000011", "0000011", "0000011", "0000101", "0000011", "0000100", "0000100", "0001010", "0000110", "0000011", "0000010", "0000110", "0001011", "0000111", "0000111", "0000100", "0001001", "0000101", "0101010", "0001001", "0001000", "0000110", "0010010", "0000110", "0000111", "0001110", "0000111", "0000100", "0000011", "0000110", "0001001", "0001001", "0011001", "0000011", "0000110", "0000011", "0000100", "0000101", "0000101", "0000010", "0000110", "0000110", "0000100", "0000101", "0000100", "0000001", "0000001", "0000101", "0010011", "0011011", "0001101", "0011000", "0100110", "0110001", "0011010", "0100111", "0010101", "0100001", "0011010", "0011100", "0100010", "0010101", "0001000", "0100101", "0100110", "0011110", "0011010", "0101100", "0011000", "0001110", "0100001", "0100011", "0010000", "0011110", "0001001", "0001100", "0001001", "0001001", "0001001", "0001001", "0001010", "0000111", "0000110", "0000111", "0000111", "0001010", "0001011", "0001111", "0000101", "0001011", "0001101", "0000011", "0011101", "0001011", "0000101", "0000011", "0001000", "0001000", "0010000", "0010001", "0001001", "0001001", "0000110", "0000111", "0000111", "0000111", "0001010", "0001101", "0001010", "0000110", "0000100", "0001110", "0011001", "0010101", "0010110", "0001011", "0010101", "0001110", "0101011", "0011000", "0010001", "0010001", "0011111", "0010001", "0010010", "0001111", "0010011", "0001011", "0000111", "0010101", "0001101", "0011010", "0011110", "0001111", "0011010", "0001010", "0010000", "0010101", "0010100", "0001001", "0011000", "0011001", "0001010", "0010000", "0001110", "0000011", "0000011", "0001101", "0010101", "0011111", "0010000", "0011100", "0100111", "0110100", "0011101", "0101110", "0010110", "0100111", "0011100", "0100000", "0101110", "0011101", "0001100", "0110101", "0111100", "0101101", "0011110", "0110100", "0011111", "0010100", "0100100", "0101011", "0010101", "0100111", "0001011", "0010010", "0001101", "0001110", "0001110", "0001111", "0010000", "0001011", "0001000", "0001101", "0001011", "0001011", "0010000", "0010101", "0000111", "0010000", "0001100", "0000101", "0100011", "0010000", "0001001", "0000101", "0001010", "0001001", "0010101", "0010010", "0001100", "0001010", "0001000", "0001001", "0001100", "0001100", "0010111", "0011010", "0010111", "0001101", "0001010", "0011010", "0001100", "0001001", "0001001", "0000101", "0001001", "0000110", "0001110", "0001100", "0001000", "0001000", "0010100", "0000111", "0001001", "0000101", "0001001", "0000101", "0000100", "0001010", "0001001", "0001011", "0001001", "0000111", "0001101", "0000101", "0001011", "0001110", "0001110", "0001011", "0011011", "0011000", "0010011", "0011101", "0011010", "0001001", "0001010", "0100100", "0001111", "0010001", "0000101", "0001010", "0001100", "0010000", "0001001", "0001101", "0001000", "0001100", "0001001", "0001010", "0001111", "0001010", "0000100", "0010110", "0011011", "0010101", "0001001", "0100110", "0011000", "0001101", "0100010", "0101000", "0010011", "0101010", "0001100", "0010011", "0011100", "0011110", "0100001", "0011111", "0100101", "0010111", "0010001", "0011000", "0010111", "0000011", "0100100", "0100100", "0010000", "0100100", "0010001", "0001100", "0001010", "0100100", "0010100", "0001010", "0011100", "0010100", "0100000", "0000110", "0100011", "0100001", "0011100", "0010000", "0100001", "0100001", "0010001", "0010111", "0010100", "0001111", "0001010", "0011111", "0000111", "0000011", "0000011", "0000001", "0000011", "0000010", "0000011", "0000011", "0000011", "0000010", "0001010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000011", "0000010", "0000101", "0000011", "0000010", "0000010", "0000100", "0000010", "0000011", "0000100", "0000100", "0000011", "0000111", "0000111", "0000110", "0001001", "0001000", "0000011", "0000011", "0001010", "0001011", "0001100", "0000001", "0000011", "0000011", "0000011", "0000010", "0000011", "0000001", "0000011", "0000010", "0000010", "0000100", "0000011", "0000001", "0000100", "0000100", "0000011", "0000010", "0000101", "0000100", "0000010", "0000111", "0001000", "0000100", "0001010", "0000101", "0000101", "0000110", "0000110", "0000110", "0000111", "0000111", "0000101", "0000100", "0000101", "0000101", "0000001", "0001000", "0001111", "0000100", "0001001", "0001011", "0000010", "0000010", "0001000", "0000100", "0000011", "0001000", "0000111", "0001111", "0000001", "0010000", "0010000", "0001100", "0001010", "0010011", "0010010", "0000010", "0000101", "0000011", "0000010", "0000010", "0000101", "0000111", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0001000", "0000000", "0000001", "0000010", "0000001", "0000000", "0000010", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000011", "0000011", "0000001", "0000001", "0000100", "0001011", "0001001", "0000000", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000010", "0000000", "0000001", "0000011", "0000010", "0000000", "0000010", "0000010", "0000001", "0000001", "0000011", "0000011", "0000001", "0000010", "0000011", "0000010", "0000011", "0000100", "0000011", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000011", "0000000", "0000010", "0001100", "0000010", "0000011", "0000111", "0000001", "0000001", "0000011", "0000001", "0000010", "0000010", "0000010", "0001001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000011", "0000011", "0000001", "0000100", "0000011", "0000001", "0000001", "0000011", "0001000", "0000010", "0000010", "0000001", "0000010", "0000010", "0000011", "0000011", "0000010", "0000010", "0001000", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000010", "0000100", "0000010", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000000", "0000001", "0001011", "0001011", "0000001", "0000011", "0000011", "0000100", "0000010", "0000011", "0000010", "0000100", "0000010", "0000011", "0000101", "0000010", "0000000", "0000010", "0000001", "0000001", "0000010", "0000001", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000010", "0001001", "0001010", "0001011", "0001011", "0001011", "0000111", "0000110", "0001000", "0001001", "0000001", "0001100", "0010000", "0000101", "0001100", "0001000", "0000100", "0000010", "0001100", "0000110", "0000100", "0000111", "0000110", "0001010", "0000010", "0000101", "0000101", "0000100", "0000010", "0000011", "0000011", "0001100", "0001111", "0001100", "0001000", "0000110", "0010000", "0001100", "0001001", "0001001", "0000101", "0001001", "0000110", "0001010", "0001011", "0001000", "0000111", "0001101", "0000111", "0001000", "0000100", "0000111", "0000101", "0000011", "0001000", "0000110", "0001010", "0000111", "0000101", "0001000", "0000011", "0000100", "0000110", "0000110", "0000010", "0000110", "0000110", "0000011", "0000101", "0000011", "0000001", "0000001", "0000010", "0001100", "0001011", "0000011", "0000110", "0001010", "0001011", "0000110", "0001010", "0000101", "0001001", "0000110", "0000111", "0001011", "0000110", "0000010", "0001001", "0001010", "0001000", "0000111", "0001001", "0000101", "0000011", "0000101", "0000110", "0000011", "0000101", "0000100", "0000011", "0001101", "0001110", "0001101", "0001111", "0001101", "0001010", "0000111", "0001100", "0001011", "0000010", "0001111", "0010100", "0000111", "0010001", "0001001", "0000110", "0000110", "0010000", "0001001", "0000101", "0001110", "0001010", "0010000", "0000100", "0010100", "0010011", "0010000", "0001010", "0010010", "0010010", "0001101", "0001111", "0001110", "0001010", "0000111", "0010101", "0001001", "0000100", "0000100", "0000010", "0000101", "0000011", "0000011", "0000110", "0000100", "0000100", "0001001", "0000011", "0000100", "0000001", "0000100", "0000011", "0000011", "0000100", "0000100", "0000101", "0000010", "0000101", "0001001", "0000011", "0000111", "0001010", "0001001", "0000110", "0010001", "0010000", "0001010", "0001111", "0001101", "0000100", "0000100", "0010001", "0001011", "0001000", "0000001", "0000011", "0000011", "0000011", "0000010", "0000011", "0000010", "0000011", "0000010", "0000010", "0000110", "0000011", "0000001", "0001000", "0001001", "0000110", "0000010", "0001100", "0000111", "0000100", "0001011", "0001101", "0000110", "0001110", "0000101", "0000111", "0000010", "0000010", "0000011", "0000011", "0000011", "0000010", "0000010", "0000010", "0000100", "0000001", "0000011", "0001100", "0000010", "0000100", "0000101", "0000001", "0000010", "0000100", "0000010", "0000010", "0000011", "0000011", "0000111", "0000001", "0000111", "0000111", "0000101", "0000110", "0001011", "0001100", "0000010", "0000100", "0000011", "0000010", "0000001", "0000100", "0000111", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000101", "0000000", "0000001", "0000001", "0000000", "0000000", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000100", "0000100", "0000100", "0000111", "0000110", "0000011", "0000011", "0001010", "0001100", "0000101", "0000000", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000011", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000011", "0000011", "0000010", "0000011", "0000011", "0000010", "0000011", "0000011", "0000011", "0000011", "0000011", "0000010", "0000010", "0000010", "0000011", "0000000", "0000011", "0001011", "0000010", "0000100", "0000100", "0000001", "0000001", "0000100", "0000010", "0000010", "0000010", "0000010", "0000101", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000010", "0000010", "0000011", "0000011", "0000001", "0000001", "0000011", "0000111", "0000001", "0000001", "0000001", "0000001", "0000001", "0000111", "0000010", "0000001", "0000000", "0000101", "0000000", "0000001", "0000011", "0000000", "0000000", "0000010", "0000001", "0000010", "0000001", "0000101", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000000", "0000001", "0001101", "0001000", "0000010", "0000101", "0000111", "0001000", "0000100", "0000110", "0000100", "0000110", "0000100", "0000101", "0000101", "0000011", "0000001", "0000010", "0000010", "0000010", "0000101", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000100", "0000100", "0000100", "0000100", "0000101", "0000011", "0000010", "0000100", "0000100", "0000010", "0000101", "0001101", "0000010", "0000101", "0000011", "0000010", "0000101", "0000101", "0000011", "0000010", "0000100", "0000011", "0000101", "0000011", "0000100", "0000101", "0000100", "0000010", "0000100", "0000100", "0000100", "0000101", "0000101", "0000011", "0000010", "0000110", "0001001", "0000100", "0000100", "0000010", "0000100", "0000011", "0001010", "0000101", "0000011", "0000011", "0000111", "0000011", "0000011", "0000100", "0000011", "0000010", "0000011", "0000100", "0000010", "0000100", "0000110", "0000001", "0000011", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000000", "0000001", "0001100", "0001001", "0000011", "0000111", "0001010", "0001101", "0000111", "0001010", "0000101", "0001001", "0000111", "0000111", "0001011", "0000111", "0000011", "0001100", "0001101", "0001010", "0000110", "0001010", "0000111", "0000100", "0000110", "0000111", "0000011", "0000100", "0000010", "0000010", "0000010", "0000010", "0000010", "0000010", "0000011", "0000010", "0000001", "0000010", "0000011", "0000011", "0000011", "0001100", "0000001", "0000011", "0000011", "0000001", "0001000", "0000011", "0000001", "0000001", "0000011", "0000010", "0000110", "0000100", "0000101", "0000100", "0000011", "0000011", "0000101", "0000101", "0000011", "0000100", "0000011", "0000010", "0000010", "0000101", "0001010", "0000110", "0000110", "0000011", "0000110", "0000100", "0000100", "0001000", "0000101", "0000101", "0001001", "0000101", "0000110", "0000001", "0000110", "0000011", "0000011", "0000110", "0000100", "0000111", "0000011", "0000100", "0001000", "0000011", "0000100", "0000110", "0000110", "0000010", "0000110", "0000110", "0000010", "0000100", "0000011", "0000001", "0000001", "0000011", "0001100", "0000101", "0000001", "0000011", "0000100", "0000101", "0000010", "0000100", "0000010", "0000011", "0000010", "0000011", "0000101", "0000010", "0000001", "0001000", "0001000", "0000110", "0000011", "0001111", "0001000", "0000100", "0001110", "0001111", "0000111", "0010000", "0000100", "0000111", "0000010", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000010", "0000010", "0000001", "0000010", "0001100", "0000001", "0000011", "0000011", "0000001", "0000011", "0000011", "0000001", "0000001", "0000001", "0000001", "0000101", "0000010", "0000010", "0000010", "0000001", "0000010", "0000011", "0000010", "0000001", "0000011", "0000011", "0000001", "0000001", "0000010", "0001001", "0000101", "0000100", "0000010", "0000100", "0000011", "0000110", "0000110", "0000011", "0000100", "0000111", "0000011", "0000100", "0000010", "0000100", "0000010", "0000011", "0000101", "0000011", "0000101", "0000100", "0000011", "0000101", "0000010", "0000100", "0000110", "0000101", "0000100", "0001011", "0001010", "0000111", "0001011", "0001001", "0000011", "0000011", "0001011", "0001011", "0000101", "0000010", "0000100", "0000101", "0000110", "0000100", "0000101", "0000011", "0000101", "0000011", "0000100", "0000101", "0000011", "0000001", "0000101", "0000101", "0000100", "0000100", "0000101", "0000011", "0000010", "0000100", "0000101", "0000010", "0000111", "0000010", "0000011", "0000101", "0000101", "0000110", "0000110", "0000111", "0000101", "0000100", "0000101", "0000101", "0000001", "0000111", "0001101", "0000011", "0001000", "0000011", "0000010", "0000100", "0000111", "0000100", "0000010", "0000100", "0000011", "0000110", "0000010", "0000100", "0000100", "0000011", "0000010", "0000010", "0000010", "0000101", "0000101", "0000101", "0000010", "0000010", "0000101", "0000101", "0000100", "0000100", "0000010", "0000100", "0000011", "0000010", "0000101", "0000011", "0000011", "0000101", "0000011", "0000011", "0000001", "0000100", "0000010", "0000010", "0000100", "0000010", "0000100", "0000001", "0000011", "0000110", "0000010", "0000100", "0000101", "0000101", "0000011", "0000110", "0000111", "0000100", "0000110", "0000110", "0000010", "0000010", "0001001", "0000100", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000011", "0000010", "0000001", "0000101", "0000101", "0000100", "0000001", "0001000", "0000100", "0000010", "0000110", "0000111", "0000011", "0000110", "0000001", "0000011", "0000011", "0000011", "0000011", "0000011", "0000011", "0000010", "0000010", "0000010", "0000010", "0000000", "0000011", "0000101", "0000010", "0000100", "0000001", "0000001", "0000001", "0000100", "0000010", "0000001", "0000100", "0000011", "0000101", "0000001", "0000111", "0000111", "0000110", "0000100", "0000111", "0000111", "0000101", "0000110", "0000110", "0000100", "0000011", "0001010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000011", "0000011", "0000011", "0000111", "0000110", "0000101", "0000111", "0000111", "0000010", "0000010", "0001000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000011", "0000100", "0000010", "0000110", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000010", "0000010", "0000010", "0000010", "0000100", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000011", "0000011", "0000001", "0000001", "0000110", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000010", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000010", "0000010", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000010", "0000001", "0000000", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000010", "0000010", "0000010", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000010", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000010", "0000010", "0000010", "0000010", "0000100", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000010", "0000011", "0000100", "0000100", "0000010", "0000010", "0000110", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000110", "0000111", "0000111", "0000100", "0000011", "0001010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000011", "0000100", "0000100", "0000011", "0001000", "0000111", "0000101", "0000111", "0000110", "0000010", "0000010", "0001000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000011", "0000010", "0000001", "0000100", "0000101", "0000010", "0000110", "0000010", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000011", "0000011", "0000010", "0000011", "0000101", "0000101", "0000100", "0000100", "0000100", "0000010", "0000001", "0000100", "0000110", "0000100", "0000100", "0000010", "0000100", "0000011", "0000010", "0000110", "0000100", "0000100", "0000110", "0000011", "0000100", "0000001", "0000100", "0000010", "0000010", "0000101", "0000010", "0000101", "0000001", "0000011", "0000110", "0000010", "0000100", "0000101", "0000100", "0000011", "0000111", "0000110", "0000101", "0001000", "0000110", "0000011", "0000011", "0001010", "0000110", "0000011", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000011", "0000010", "0000001", "0000110", "0000110", "0000101", "0000001", "0001000", "0000100", "0000010", "0000101", "0000111", "0000011", "0000101", "0000001", "0000010", "0000100", "0000100", "0000100", "0000100", "0000101", "0000011", "0000011", "0000100", "0000011", "0000001", "0000101", "0001000", "0000010", "0000101", "0000010", "0000010", "0000010", "0000101", "0000011", "0000001", "0000101", "0000011", "0000110", "0000001", "0001000", "0000111", "0000110", "0000100", "0000110", "0000110", "0000001", "0000011", "0000011", "0000001", "0000001", "0000010", "0001000", "0000100", "0000100", "0000010", "0000100", "0000011", "0000110", "0000101", "0000011", "0000100", "0000111", "0000011", "0000100", "0000010", "0000100", "0000010", "0000011", "0000100", "0000011", "0000101", "0000100", "0000011", "0000110", "0000010", "0000101", "0000111", "0000110", "0000100", "0001011", "0001011", "0000110", "0001010", "0001001", "0000010", "0000011", "0001001", "0001100", "0000101", "0000010", "0000100", "0000101", "0000111", "0000100", "0000110", "0000011", "0000101", "0000100", "0000100", "0000101", "0000011", "0000001", "0000100", "0000101", "0000100", "0000100", "0000101", "0000011", "0000010", "0000110", "0000110", "0000011", "0001001", "0000011", "0000100", "0000101", "0000101", "0000110", "0000101", "0000110", "0000100", "0000011", "0000101", "0000100", "0000001", "0000110", "0001101", "0000011", "0000111", "0000100", "0000010", "0000100", "0000110", "0000011", "0000010", "0000011", "0000011", "0000101", "0000011", "0000011", "0000011", "0000010", "0000001", "0000010", "0000010", "0000011", "0000100", "0000100", "0000011", "0000010", "0000101", "0001010", "0000111", "0000111", "0000100", "0000111", "0000101", "0000100", "0001000", "0000110", "0000101", "0001001", "0000101", "0000110", "0000010", "0000110", "0000011", "0000011", "0000111", "0000100", "0001000", "0000011", "0000100", "0000111", "0000011", "0000100", "0000101", "0000101", "0000010", "0000101", "0000100", "0000010", "0000011", "0000010", "0000000", "0000001", "0000010", "0001011", "0000110", "0000001", "0000011", "0000100", "0000101", "0000011", "0000100", "0000010", "0000011", "0000011", "0000011", "0000101", "0000011", "0000001", "0001001", "0001011", "0001000", "0000010", "0010000", "0001010", "0000101", "0001110", "0010000", "0000111", "0001111", "0000100", "0000110", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0001100", "0000001", "0000010", "0000011", "0000001", "0000011", "0000011", "0000001", "0000001", "0000001", "0000001", "0000110", "0000010", "0000010", "0000010", "0000010", "0000010", "0000011", "0000011", "0000100", "0000101", "0000101", "0000010", "0000010", "0000101", "0001000", "0000011", "0000011", "0000010", "0000011", "0000010", "0001011", "0000100", "0000010", "0000010", "0000110", "0000010", "0000011", "0000100", "0000010", "0000001", "0000011", "0000011", "0000010", "0000011", "0001000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0001101", "0001001", "0000100", "0001000", "0001011", "0001110", "0000111", "0001011", "0000110", "0001010", "0001000", "0001000", "0001011", "0000110", "0000011", "0001011", "0001011", "0001000", "0000111", "0001000", "0000101", "0000011", "0000011", "0000100", "0000010", "0000010", "0000010", "0000010", "0000011", "0000011", "0000011", "0000011", "0000011", "0000010", "0000010", "0000010", "0000011", "0000011", "0000011", "0001100", "0000010", "0000100", "0000011", "0000001", "0001001", "0000100", "0000010", "0000001", "0000011", "0000010", "0000110", "0000101", "0000101", "0000101", "0000011", "0000011", "0000101", "0000101", "0000010", "0000011", "0000011", "0000001", "0000001", "0000011", "0000111", "0000001", "0000000", "0000000", "0000001", "0000001", "0000101", "0000010", "0000001", "0000000", "0000101", "0000000", "0000001", "0000010", "0000000", "0000000", "0000010", "0000001", "0000010", "0000001", "0000011", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000000", "0000001", "0001100", "0000111", "0000010", "0000100", "0000101", "0000110", "0000011", "0000101", "0000010", "0000100", "0000011", "0000100", "0000100", "0000010", "0000001", "0000010", "0000010", "0000001", "0000011", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000100", "0000100", "0000100", "0000100", "0000101", "0000011", "0000010", "0000100", "0000100", "0000001", "0000101", "0001101", "0000010", "0000101", "0000011", "0000010", "0000100", "0000101", "0000011", "0000010", "0000100", "0000011", "0000101", "0000010", "0000100", "0000100", "0000011", "0000010", "0000011", "0000011", "0000011", "0000101", "0000100", "0000011", "0000010", "0000111", "0000111", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000101", "0000000", "0000001", "0000001", "0000001", "0000000", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000011", "0000110", "0000110", "0000110", "0001011", "0001000", "0000011", "0000100", "0001110", "0001100", "0000101", "0000000", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000100", "0000001", "0000000", "0000010", "0000010", "0000001", "0000001", "0000100", "0000010", "0000001", "0000100", "0000110", "0000011", "0000110", "0000011", "0000100", "0000010", "0000011", "0000011", "0000010", "0000011", "0000010", "0000010", "0000010", "0000011", "0000000", "0000011", "0001011", "0000010", "0000100", "0000100", "0000001", "0000001", "0000100", "0000010", "0000010", "0000010", "0000010", "0000110", "0000000", "0000010", "0000010", "0000010", "0000010", "0000010", "0000011", "0001111", "0010001", "0001111", "0001011", "0001000", "0011000", "0001010", "0000110", "0000110", "0000011", "0000110", "0000100", "0000100", "0001001", "0000110", "0000101", "0001011", "0000100", "0000110", "0000010", "0000110", "0000011", "0000011", "0000110", "0000101", "0001000", "0000011", "0000110", "0001010", "0000100", "0001000", "0001011", "0001010", "0000110", "0010000", "0010000", "0001000", "0001101", "0001100", "0000100", "0000100", "0001101", "0001011", "0001001", "0000001", "0000100", "0000100", "0000101", "0000011", "0000100", "0000010", "0000100", "0000011", "0000011", "0001000", "0000100", "0000001", "0001001", "0001011", "0001000", "0000011", "0001101", "0001000", "0000101", "0001100", "0001101", "0000110", "0001101", "0000101", "0000110", "0000011", "0000011", "0000011", "0000011", "0000100", "0000010", "0000010", "0000011", "0000100", "0000001", "0000100", "0001101", "0000011", "0000101", "0000110", "0000001", "0000011", "0000101", "0000010", "0000010", "0000101", "0000100", "0001000", "0000010", "0001010", "0001010", "0001000", "0000111", "0001110", "0001110", "0001001", "0001100", "0001010", "0000101", "0000011", "0001010", "0001011", "0000111", "0001000", "0000100", "0001000", "0000101", "0001010", "0001001", "0000110", "0000110", "0001011", "0000110", "0000111", "0000100", "0000110", "0000100", "0000011", "0000111", "0000101", "0001000", "0000111", "0000011", "0000111", "0000011", "0000011", "0000100", "0000100", "0000010", "0000100", "0000100", "0000010", "0000100", "0000010", "0000000", "0000001", "0000010", "0001100", "0001011", "0000011", "0000110", "0001001", "0001011", "0000110", "0001010", "0000101", "0001000", "0000110", "0000111", "0001001", "0000101", "0000010", "0000111", "0001000", "0000110", "0000111", "0000110", "0000100", "0000010", "0000011", "0000011", "0000010", "0000011", "0000100", "0000010", "0001111", "0001111", "0010000", "0010010", "0010000", "0001011", "0001001", "0001101", "0001101", "0000011", "0010010", "0010101", "0001000", "0010010", "0001010", "0000110", "0000111", "0010011", "0001010", "0000101", "0001110", "0001011", "0010000", "0000100", "0010010", "0010010", "0001110", "0001000", "0001111", "0001111", "0000001", "0000100", "0000010", "0000001", "0000001", "0000011", "0000111", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000011", "0000010", "0000001", "0001000", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000100", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000000", "0000001", "0001011", "0001011", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000011", "0000001", "0000010", "0000100", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000010", "0000110", "0000111", "0001000", "0000111", "0000111", "0000110", "0000100", "0000110", "0000110", "0000001", "0001000", "0001110", "0000100", "0001010", "0000111", "0000011", "0000001", "0001000", "0000101", "0000011", "0000100", "0000100", "0001001", "0000001", "0000100", "0000011", "0000010", "0000010", "0000010", "0000010", "0000100", "0000111", "0000101", "0000101", "0000011", "0001010", "0000111", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000011", "0000010", "0000001", "0001000", "0000001", "0000001", "0000010", "0000001", "0000000", "0000010", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000011", "0000011", "0000010", "0000100", "0000011", "0000001", "0000001", "0000100", "0001011", "0001001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000011", "0000010", "0000000", "0000011", "0000011", "0000010", "0000001", "0000011", "0000011", "0000010", "0000011", "0000011", "0000010", "0000011", "0000100", "0000011", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000011", "0000000", "0000010", "0001100", "0000010", "0000011", "0001000", "0000001", "0000001", "0000011", "0000001", "0000010", "0000010", "0000011", "0001010", "0000001", "0000011", "0000011", "0000010", "0000010", "0000011", "0000011", "0011011", "0100000", "0011101", "0010100", "0001110", "0101010", "0001000", "0000011", "0000011", "0000010", "0000100", "0000010", "0000011", "0000101", "0000011", "0000011", "0001011", "0000011", "0000011", "0000010", "0000011", "0000010", "0000011", "0000011", "0000110", "0000100", "0000010", "0000011", "0000101", "0000010", "0000100", "0000101", "0000101", "0000100", "0001010", "0001010", "0000110", "0001010", "0001000", "0000011", "0000100", "0001110", "0001100", "0001100", "0000001", "0000011", "0000011", "0000011", "0000010", "0000011", "0000010", "0000100", "0000010", "0000010", "0000100", "0000011", "0000001", "0000100", "0000101", "0000100", "0000010", "0001001", "0000111", "0000100", "0001000", "0001011", "0000101", "0001100", "0000101", "0000110", "0001001", "0001001", "0001011", "0001011", "0001100", "0001000", "0000110", "0001000", "0001001", "0000001", "0001011", "0010001", "0000110", "0001101", "0001101", "0000100", "0000010", "0001100", "0000111", "0000100", "0001101", "0001001", "0010011", "0000001", "0010111", "0010110", "0010001", "0001101", "0011011", "0011011", "0001111", "0010010", "0010000", "0000111", "0000110", "0010000", "0010000", "0001011", "0001100", "0000110", "0001011", "0001000", "0010010", "0001111", "0001010", "0001010", "0010111", "0001001", "0001010", "0000111", "0001011", "0000110", "0000101", "0001011", "0001001", "0001110", "0001110", "0001001", "0010001", "0000110", "0001110", "0010100", "0010001", "0001100", "0011111", "0011101", "0010011", "0011101", "0011010", "0001001", "0001001", "0100010", "0010001", "0010100", "0000111", "0001100", "0010010", "0010111", "0001101", "0010100", "0001001", "0010001", "0001100", "0001101", "0010101", "0001111", "0000110", "0100010", "0101001", "0011110", "0001101", "0101011", "0011010", "0001111", "0100001", "0101000", "0010011", "0101001", "0001100", "0010011", "0011101", "0011111", "0100000", "0100000", "0100101", "0010111", "0010001", "0011001", "0010111", "0000101", "0100101", "0100111", "0001111", "0100110", "0010001", "0001011", "0001111", "0100011", "0010011", "0001001", "0011001", "0010100", "0011111", "0001000", "0011110", "0011100", "0010111", "0001111", "0011100", "0011010", "0000111", "0001011", "0000111", "0000101", "0000011", "0001001", "0010111", "0010101", "0010101", "0001011", "0010101", "0001110", "0101111", "0011000", "0010000", "0010001", "0011101", "0010000", "0010011", "0010000", "0010011", "0001011", "0000111", "0010100", "0001101", "0011001", "0011100", "0001100", "0010110", "0001000", "0001100", "0001111", "0010001", "0000111", "0010010", "0010001", "0001001", "0001110", "0001101", "0000010", "0000011", "0001011", "0010110", "0011111", "0010000", "0011110", "0101001", "0110111", "0011111", "0101101", "0011001", "0101000", "0011111", "0100001", "0101101", "0011100", "0001011", "0101100", "0110000", "0101000", "0011110", "0110001", "0011100", "0010010", "0100101", "0101011", "0010101", "0100110", "0001010", "0010001", "0001011", "0001100", "0001100", "0001100", "0001110", "0001001", "0000111", "0001001", "0001000", "0001100", "0001101", "0010000", "0000110", "0001110", "0001100", "0000100", "0100011", "0001110", "0000111", "0000100", "0001001", "0001001", "0010011", "0010100", "0001101", "0001011", "0001000", "0001000", "0001001", "0001010", "0000100", "0001001", "0000110", "0000010", "0000010", "0000110", "0001001", "0000101", "0000110", "0000011", "0000111", "0000100", "0100111", "0000111", "0000110", "0000101", "0010001", "0000100", "0000101", "0001101", "0000100", "0000011", "0000011", "0000101", "0001000", "0000111", "0011000", "0000011", "0000101", "0000010", "0000100", "0000100", "0000100", "0000010", "0000101", "0000101", "0000100", "0000101", "0000100", "0000001", "0000001", "0000110", "0010010", "0011001", "0001101", "0010111", "0100011", "0101101", "0010110", "0100101", "0010100", "0100000", "0010110", "0011011", "0100010", "0010101", "0001000", "0101000", "0101100", "0100001", "0011001", "0110000", "0011101", "0010000", "0100110", "0101001", "0010011", "0100100", "0001010", "0001111", "0001000", "0001000", "0001000", "0001001", "0001010", "0000110", "0000101", "0000111", "0000111", "0001001", "0001001", "0001111", "0000101", "0001010", "0001100", "0000011", "0011100", "0001010", "0000110", "0000011", "0000111", "0000111", "0010001", "0010000", "0000110", "0000111", "0000101", "0000110", "0000111", "0000111", "0000010", "0001001", "0000011", "0000011", "0000011", "0000111", "0001110", "0001010", "0001010", "0000110", "0001100", "0001000", "0110101", "0001101", "0001011", "0001001", "0011100", "0001000", "0001010", "0010011", "0001001", "0000101", "0000100", "0001000", "0001010", "0001011", "0100100", "0000110", "0001010", "0000100", "0001010", "0001101", "0001101", "0001001", "0011000", "0010110", "0001001", "0001101", "0001100", "0001000", "0001000", "0011111", "0011010", "0100110", "0010010", "0100010", "0110000", "0111110", "0100001", "0110101", "0011001", "0101010", "0100000", "0100011", "0101111", "0100000", "0001100", "1000000", "1000111", "0110110", "0100010", "1001001", "0101010", "0011001", "0110010", "0111100", "0011100", "1000000", "0010010", "0011101", "0000011", "0000011", "0000011", "0000011", "0000100", "0000010", "0000011", "0000011", "0000011", "0001101", "0000101", "0001100", "0000100", "0000100", "0001101", "0000001", "0101000", "0000101", "0000011", "0000011", "0000100", "0000101", "0010101", "0010110", "0000011", "0000011", "0000011", "0000110", "0000111", "0000111", "0011110", "0101010", "0100000", "0001111", "0001011", "0100010", "0101111", "0101101", "0101011", "0010110", "0101100", "0011101", "0101011", "0110011", "0100100", "0100101", "1000001", "0100001", "0101000", "0010001", "0101000", "0010110", "0001111", "0100111", "0011010", "0101110", "0100000", "0011011", "0110000", "0010010", "0100000", "0101010", "0101001", "0010011", "0110010", "0110001", "0101000", "0111011", "0110110", "0001100", "0001101", "0101111", "0010010", "0110001", "0001111", "0011101", "0101000", "0110101", "0011101", "0101010", "0011001", "0101000", "0011101", "0100001", "0101011", "0011110", "0001010", "0100011", "0100011", "0011011", "0011110", "0110000", "0011101", "0010000", "0011111", "0100010", "0010010", "0011111", "0001010", "0001101", "0011010", "0011101", "0011111", "0011110", "0100010", "0010111", "0010001", "0011000", "0010110", "0001011", "0011100", "0100001", "0001110", "0011111", "0011010", "0001011", "0100010", "0011101", "0010000", "0001000", "0010100", "0010010", "0101010", "0010100", "0100011", "0100010", "0011011", "0010001", "0011000", "0011010", "0100011", "0110100", "0100010", "0011000", "0010001", "0101111", "0100101", "0100010", "0100001", "0010010", "0100001", "0011000", "0100110", "0101010", "0011101", "0011101", "1000001", "0011010", "0011111", "0010000", "0011101", "0010001", "0001011", "0011111", "0100101", "0100110", "0011011", "0010110", "0100111", "0001110", "0010101", "0011100", "0011011", "0010011", "0110100", "0110000", "0011010", "0101000", "0100100", "0001001", "0001010", "0100101", "0010000", "0111101", "0001110", "0011001", "0100011", "0101101", "0011011", "0100111", "0010010", "0100010", "0010111", "0011100", "0011111", "0010111", "0000111", "0101011", "0110000", "0100011", "0011011", "0100101", "0011101", "0010000", "0101000", "0110010", "0011000", "0011011", "0001011", "0001101", "0101100", "0101111", "0110010", "0110100", "0110110", "0100101", "0011110", "0101010", "0100101", "0001010", "0111011", "0111001", "0011001", "0111010", "0111001", "0010010", "0011101", "0110011", "0011011", "0001101", "0101010", "0011110", "1000101", "0010001", "0101100", "0101000", "0011111", "0100000", "0110101", "0110100", "0001010", "0000000", "0000101", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0001111", "0000101", "0001010", "0000101", "0000101", "0000000", "0000101", "0000101", "0001010", "0000101", "0011001", "0000000", "0000000", "0010100", "0001010", "0001010", "0001111", "0000101", "0000101", "0001010", "0001010", "0001010", "0000000", "0000101", "0000101", "0001111", "0001010", "0000000", "0000101", "0000000", "0000000", "0000101", "0001010", "0001010", "0000101", "0000101", "0001111", "0000000", "0001010", "0001111", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000101", "0001010", "0001010", "0000101", "0000000", "0001010", "0001010", "0001010", "0001010", "0001010", "0001010", "0010100", "0000101", "0001111", "0001010", "0000000", "0001010", "0001010", "0000000", "0000101", "0000101", "0001111", "0001111", "0000101", "0000000", "0001111", "0100011", "0011001", "0000101", "0011001", "0000000", "0001111", "0001010", "0000101", "0000101", "0000000", "0000000", "0010100", "0000000", "0100011", "0010001", "0101100", "0010010", "0010111", "0011100", "0001100", "0010010", "0001100", "0011100", "0010110", "0110011", "0010010", "0100101", "0010101", "0101010", "0001101", "0100011", "0011010", "1000010", "0001111", "0010111", "0111101", "0101010", "0111000", "0010100", "0011100", "0010001", "0100010", "0011000", "0010011", "0001010", "0001010", "0011110", "0100111", "0011110", "0001011", "0011011", "0001100", "0010101", "0011001", "0010011", "0010111", "0001100", "0010000", "0100000", "0001001", "0011000", "0100010", "0001000", "0101011", "0001101", "0010000", "0001010", "0010011", "0001101", "0011111", "0100000", "0011000", "0011011", "0001110", "0010110", "0110011", "0101101", "0010001", "0011100", "0010011", "0100010", "0011110", "0100010", "0101101", "0101110", "0110010", "0011000", "0100110", "0001111", "0010000", "0101100", "0011110", "0010110", "0110001", "0011101", "0101011", "0110101", "0100011", "0011000", "1010001", "1001001", "0110010", "0010010", "0110001", "0001011", "0101100", "0110100", "0010100", "0101100", "0011010", "0011101", "1001100", "0100000", "0011010", "0101001", "1001111", "0100111", "0110101", "1011110", "0100000", "0111100", "0100110", "0100000", "0001110", "0100001", "0001011", "0010110", "0001101", "0011001", "0001001", "0010100", "0011111", "0101000", "0001001", "0010001", "0111011", "0011100", "0100000", "0010001", "0011111", "0010011", "0100101", "0010011", "0010100", "0001010", "0001100", "0100011", "0101000", "0100010", "0001101", "0100001", "0001101", "0010111", "0011010", "0010101", "0011001", "0001110", "0010010", "0100110", "0001011", "0011101", "0100111", "0001001", "0100101", "0001011", "0001110", "0001001", "0011000", "0001111", "0100110", "0100110", "0011110", "0100000", "0001111", "0011000", "0110100", "0110000", "0010010", "0011101", "0010101", "0100101", "0100001", "0011011", "0101010", "0110010", "0110100", "0011010", "0101010", "0010000", "0010001", "0101111", "0011111", "0010111", "0110100", "0100001", "0101101", "0111101", "0100110", "0011001", "1001110", "1010110", "0111110", "0010111", "0111111", "0001011", "1000111", "1010111", "0100010", "0101010", "0011110", "0100000", "1001110", "0100110", "0010111", "0000010", "0001000", "0000100", "0000011", "0001001", "0000100", "0000110", "0000100", "0011100", "0000100", "0000101", "0000011", "0000010", "0000001", "0000010", "0000010", "0000001", "0011010", "0000010", "0000010", "0000110", "0100100", "0001000", "0000011", "0001111", "0011010", "0010001", "0100001", "0010001", "0010010", "0001001", "0001010", "0011101", "0011010", "0011101", "0001011", "0011100", "0001011", "0010011", "0010101", "0010011", "0010110", "0001101", "0010000", "0011111", "0001001", "0010111", "0100000", "0000111", "0110100", "0001111", "0010011", "0001100", "0010011", "0001100", "0011111", "0011111", "0101100", "0101110", "0001111", "0011100", "0000011", "0000011", "0000010", "0000010", "0010010", "0000011", "0000010", "0000111", "0011010", "0000110", "0000011", "0000011", "0000011", "0001101", "0000010", "0000011", "0000011", "0000010", "0000011", "0000110", "0011110", "0010001", "0001000", "0000010", "0101000", "0010000", "0000100", "0000001", "0000101", "0001010", "0000100", "0000100", "0000010", "0010101", "0000011", "0000100", "0100111", "0000011", "0001010", "0000000", "0000101", "0000011", "0000001", "0000001", "0000010", "0000001", "0000001", "0000100", "0000011", "0000100", "0000010", "0000001", "0000000", "0000001", "0000010", "0000001", "0000011", "0000001", "0000001", "0000100", "0010110", "0000101", "0000001", "0000100", "0000100", "0000010", "0000101", "0000101", "0000100", "0000010", "0000010", "0000100", "0001101", "0000100", "0000001", "0000011", "0000010", "0000100", "0000101", "0000011", "0000100", "0000010", "0000011", "0001000", "0000010", "0000101", "0000111", "0000001", "0000110", "0000010", "0000010", "0000010", "0000101", "0000100", "0001000", "0001000", "0001010", "0001110", "0000110", "0001001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000010", "0000001", "0000110", "0001110", "0000100", "0000001", "0000010", "0000001", "0000110", "0000001", "0000001", "0000001", "0000010", "0000001", "0000100", "0010000", "0001100", "0000100", "0000001", "0010100", "0000111", "0000001", "0000000", "0000011", "0000011", "0000001", "0000001", "0000000", "0001100", "0000001", "0000010", "0010101", "0000001", "0000110", "0000000", "0000100", "0000010", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000010", "0000011", "0000010", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000100", "0010100", "0000101", "0000001", "0000010", "0000001", "0000000", "0000001", "0000011", "0000011", "0000010", "0000001", "0000010", "0001101", "0000001", "0000000", "0000001", "0000001", "0000010", "0000011", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000111", "0000100", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000100", "0001011", "0000100", "0000001", "0000010", "0000001", "0000110", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0001111", "0001001", "0000011", "0000001", "0010001", "0000110", "0000001", "0000000", "0000011", "0000100", "0000001", "0000001", "0000000", "0001011", "0000001", "0000010", "0010110", "0000000", "0000100", "0000000", "0000011", "0000010", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000011", "0010110", "0000110", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000011", "0000001", "0000001", "0000010", "0001110", "0000001", "0000000", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000111", "0000011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0001100", "0000011", "0000001", "0000010", "0000001", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0001111", "0001011", "0000011", "0000001", "0010011", "0000111", "0000001", "0000000", "0000010", "0000011", "0000001", "0000001", "0000000", "0001011", "0000000", "0000010", "0011011", "0000000", "0000101", "0000000", "0000010", "0000010", "0000001", "0000000", "0000010", "0000000", "0000000", "0000110", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000101", "0000001", "0000001", "0000011", "0010011", "0000011", "0000001", "0000100", "0000110", "0000011", "0000111", "0000100", "0000101", "0000011", "0000010", "0000110", "0001100", "0000111", "0000010", "0000110", "0000010", "0000100", "0000101", "0000010", "0000011", "0000001", "0000010", "0000011", "0000001", "0000010", "0000011", "0000010", "0000011", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000111", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000010", "0001010", "0000010", "0000001", "0000010", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0001010", "0001000", "0000011", "0000000", "0010000", "0000110", "0000001", "0000000", "0000010", "0000010", "0000000", "0000001", "0000000", "0001001", "0000000", "0000010", "0001111", "0000000", "0010010", "0000001", "0000010", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0011001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0011000", "0000001", "0000010", "0000011", "0001100", "0000010", "0000001", "0001110", "0011001", "0001111", "0011110", "0001111", "0010000", "0000111", "0001001", "0011010", "0001011", "0011010", "0001010", "0010111", "0001010", "0010000", "0010010", "0001111", "0010010", "0001010", "0001101", "0010111", "0000110", "0010001", "0011000", "0000111", "0011001", "0000111", "0001001", "0000110", "0001001", "0000110", "0010000", "0010000", "0001110", "0010000", "0000101", "0001001", "0000101", "0000101", "0000010", "0000011", "0001111", "0000100", "0000011", "0000100", "0001001", "0000101", "0000101", "0000100", "0000100", "0001001", "0000010", "0000100", "0000011", "0000011", "0000101", "0000100", "0010001", "0001001", "0000100", "0000010", "0001111", "0000111", "0000011", "0000001", "0000100", "0000111", "0000010", "0000010", "0000001", "0000111", "0000001", "0000011", "0001101", "0000001", "0001011", "0000111", "0001100", "0000111", "0001000", "0001011", "0000100", "0000111", "0000100", "0001111", "0000101", "0001011", "0000100", "0001000", "0000101", "0001001", "0000100", "0001000", "0001101", "0001110", "0000100", "0000110", "0001101", "0001000", "0001011", "0000111", "0001101", "0001001", "0010001", "0001000", "0001010", "0000100", "0000101", "0001111", "0001000", "0001111", "0000110", "0001110", "0000110", "0001001", "0001010", "0001011", "0001100", "0000111", "0001001", "0010111", "0000111", "0010001", "0011000", "0000100", "0100100", "0001011", "0001101", "0001000", "0010101", "0001100", "0100000", "0100001", "0100110", "0101000", "0001100", "0010111", "0011100", "0011001", "0001010", "0001111", "0001001", "0010010", "0010001", "0001110", "0001001", "0011001", "0011011", "0001110", "0010101", "0000110", "0001000", "0010111", "0010000", "0001100", "0011011", "0010000", "0001010", "0011100", "0010010", "0001101", "0010110", "0100110", "0011100", "0001010", "0011101", "0000101", "0010111", "0011110", "0001011", "0001001", "0001000", "0001011", "0010001", "0001011", "0000110", "0010001", "0011110", "0010000", "0010101", "0101100", "0001111", "0011011", "0010001", "0001000", "0001010", "0011001", "0001000", "0010010", "0001011", "0010101", "0000111", "0010001", "0001000", "0100000", "0000111", "0001011", "0010001", "0010011", "0011011", "0000100", "0001000", "0000101", "0001010", "0000101", "0000101", "0000010", "0000011", "0001001", "0000101", "0001000", "0000011", "0001000", "0000011", "0000110", "0000110", "0000110", "0000111", "0000100", "0000101", "0001011", "0000011", "0001001", "0001011", "0000010", "0010001", "0000101", "0000110", "0000100", "0001001", "0000111", "0010000", "0001111", "0010001", "0010001", "0000110", "0001010", "0000111", "0000110", "0000010", "0000100", "0000110", "0000101", "0000100", "0000100", "0000110", "0000110", "0000111", "0000100", "0000101", "0000011", "0000010", "0000110", "0000100", "0000100", "0000111", "0000100", "0001000", "0001000", "0000101", "0000011", "0001011", "0010000", "0001011", "0000100", "0001011", "0000011", "0010001", "0010011", "0000111", "0001000", "0001100", "0001101", "0010101", "0001110", "0001010", "0000011", "0000101", "0000101", "0000011", "0000111", "0000101", "0000101", "0000011", "0001110", "0000011", "0001001", "0000010", "0000110", "0000100", "0000111", "0000100", "0000101", "0001110", "0001010", "0000100", "0000101", "0001011", "0000110", "0001000", "0001000", "0001110", "0001001", "0010001", "0001001", "0001001", "0000100", "0000101", "0001111", "0001000", "0010000", "0000110", "0001110", "0000110", "0001010", "0001011", "0001000", "0001001", "0000101", "0000111", "0001010", "0000011", "0001001", "0001100", "0000100", "0001100", "0000100", "0000100", "0000011", "0000110", "0000101", "0001011", "0001010", "0001100", "0001110", "0000100", "0001000", "0001111", "0001110", "0000101", "0001001", "0001010", "0001010", "0001001", "0001000", "0001000", "0001110", "0010000", "0001000", "0001100", "0000101", "0000101", "0001110", "0001001", "0000111", "0001111", "0001001", "0001011", "0001110", "0001010", "0000111", "0010000", "0001110", "0001011", "0000100", "0001011", "0000101", "0000110", "0000111", "0000011", "0000110", "0000010", "0000110", "0001011", "0000011", "0001001", "0001010", "0010011", "0001011", "0001101", "0010001", "0000110", "0001011", "0000111", "0001101", "0000111", "0010011", "0000110", "0001110", "0001000", "0001111", "0000101", "0001101", "0001100", "0011000", "0000110", "0001001", "0001110", "0001110", "0010100", "0000111", "0001011", "0000111", "0001101", "0000111", "0001000", "0000011", "0000101", "0001101", "0000110", "0001101", "0000101", "0001011", "0000101", "0001000", "0001001", "0001001", "0001011", "0000110", "0001000", "0010011", "0000101", "0001110", "0010010", "0000011", "0011010", "0001000", "0001001", "0000110", "0001101", "0001000", "0010101", "0010101", "0010101", "0010101", "0000110", "0001101", "0010110", "0010100", "0000111", "0001011", "0001000", "0001111", "0001110", "0001011", "0001000", "0010100", "0010110", "0001011", "0010001", "0000101", "0000110", "0010010", "0001100", "0001001", "0010100", "0001100", "0001001", "0010111", "0001111", "0001010", "0010010", "0100110", "0011100", "0001011", "0011100", "0000100", "0011110", "0100001", "0001110", "0001010", "0001100", "0001111", "0010100", "0001111", "0000011", "0001110", "0011100", "0001110", "0010001", "0101000", "0001110", "0011001", "0010000", "0000100", "0000011", "0000110", "0000010", "0000100", "0000011", "0000101", "0000011", "0000100", "0000100", "0001001", "0000011", "0000100", "0001001", "0000101", "0000111", "0000010", "0000100", "0000011", "0000101", "0000011", "0000011", "0000001", "0000001", "0000101", "0000101", "0000100", "0000010", "0000100", "0000010", "0000010", "0000011", "0000100", "0000101", "0000011", "0000100", "0001010", "0000011", "0000111", "0001011", "0000001", "0010010", "0000101", "0000110", "0000100", "0001010", "0000111", "0010000", "0010000", "0010100", "0010101", "0000111", "0001100", "0000010", "0000010", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000100", "0000010", "0000010", "0000011", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000010", "0000010", "0000101", "0000100", "0000010", "0000001", "0000111", "0001000", "0000101", "0000010", "0000101", "0000001", "0001001", "0001100", "0000100", "0000101", "0001001", "0001001", "0001101", "0001011", "0000001", "0000001", "0000011", "0000011", "0000010", "0000110", "0000011", "0000011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000110", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000011", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000000", "0000010", "0000010", "0000000", "0000100", "0000001", "0000010", "0000001", "0000011", "0000011", "0000111", "0000110", "0001010", "0001101", "0000011", "0000111", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000011", "0000010", "0000001", "0000110", "0000010", "0000010", "0000000", "0000010", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000010", "0000110", "0000001", "0000100", "0000000", "0000001", "0000011", "0000001", "0000001", "0000010", "0000001", "0000001", "0000101", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000101", "0000001", "0000001", "0000001", "0000110", "0000001", "0000001", "0000011", "0000101", "0000011", "0000111", "0000011", "0000100", "0000010", "0000010", "0000110", "0000100", "0000110", "0000010", "0000101", "0000010", "0000100", "0000101", "0000010", "0000010", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000010", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000001", "0001011", "0001011", "0000100", "0000111", "0000100", "0001000", "0000111", "0000110", "0000100", "0001010", "0001011", "0000110", "0001001", "0000010", "0000100", "0001010", "0000110", "0000101", "0001010", "0000110", "0000101", "0001011", "0000111", "0000101", "0001010", "0001000", "0000110", "0000010", "0000110", "0000010", "0000010", "0000011", "0000001", "0000011", "0000001", "0000010", "0000110", "0000001", "0000111", "0000100", "0000111", "0000100", "0000101", "0000100", "0000010", "0000011", "0000010", "0001010", "0000011", "0001000", "0000011", "0000111", "0000011", "0000111", "0000010", "0000110", "0001001", "0001010", "0000010", "0000100", "0001000", "0000110", "0001000", "0000101", "0001010", "0000110", "0001100", "0000110", "0000111", "0000011", "0000011", "0001010", "0000100", "0001010", "0000100", "0001010", "0000100", "0000111", "0000111", "0000111", "0001000", "0000101", "0000110", "0001010", "0000011", "0001000", "0001011", "0000011", "0001001", "0000010", "0000011", "0000010", "0000010", "0000010", "0000100", "0000100", "0000010", "0000111", "0000001", "0000010", "0010001", "0001111", "0000110", "0001001", "0000110", "0001011", "0001011", "0001000", "0000101", "0001111", "0010001", "0001001", "0001101", "0000100", "0000101", "0001111", "0001010", "0000111", "0010000", "0001001", "0000111", "0010001", "0001011", "0001000", "0001101", "0011100", "0010100", "0000111", "0010100", "0000011", "0010010", "0010110", "0001001", "0000110", "0000111", "0000111", "0001011", "0001000", "0000101", "0001100", "0010111", "0001100", "0010000", "0011100", "0001001", "0010000", "0001011", "0000111", "0000100", "0001001", "0000011", "0000111", "0000100", "0001000", "0000010", "0000111", "0000111", "0001101", "0000011", "0000100", "0000111", "0001000", "0001011", "0000100", "0000111", "0000100", "0001000", "0000100", "0000101", "0000010", "0000011", "0001000", "0000011", "0001000", "0000011", "0000111", "0000011", "0000101", "0000110", "0000101", "0000101", "0000011", "0000100", "0001010", "0000011", "0000111", "0001010", "0000010", "0001111", "0000101", "0000110", "0000100", "0001001", "0000101", "0001110", "0001110", "0001111", "0010000", "0000100", "0001001", "0001110", "0001100", "0000100", "0000111", "0000101", "0001001", "0001000", "0000111", "0000101", "0001100", "0001101", "0000110", "0001011", "0000011", "0000100", "0001011", "0000111", "0000101", "0001101", "0000111", "0000110", "0001101", "0001001", "0000110", "0001011", "0010011", "0001110", "0000101", "0001101", "0000010", "0001111", "0010010", "0000111", "0000101", "0001001", "0001010", "0001110", "0001100", "0000011", "0000111", "0001110", "0000110", "0001001", "0010001", "0000110", "0001100", "0000111", "0000100", "0000100", "0001010", "0000011", "0000110", "0000100", "0001000", "0000010", "0000110", "0000100", "0001100", "0000011", "0000100", "0000110", "0000111", "0001001", "0000010", "0000100", "0000011", "0000101", "0000010", "0000011", "0000001", "0000001", "0000100", "0000010", "0000100", "0000010", "0000100", "0000010", "0000011", "0000011", "0000100", "0000101", "0000011", "0000011", "0001001", "0000010", "0000110", "0001001", "0000001", "0001011", "0000011", "0000100", "0000011", "0000110", "0000011", "0001001", "0001001", "0001011", "0001011", "0000011", "0000111", "0000101", "0000100", "0000010", "0000011", "0000011", "0000100", "0000011", "0000011", "0000010", "0000101", "0000101", "0000011", "0000100", "0000001", "0000010", "0000101", "0000011", "0000010", "0000101", "0000011", "0000011", "0000110", "0000100", "0000011", "0000101", "0001111", "0001010", "0000100", "0001010", "0000001", "0001110", "0010001", "0000110", "0000100", "0000111", "0001000", "0001011", "0001001", "0000001", "0000111", "0001100", "0000111", "0001000", "0010011", "0000110", "0001100", "0000111", "0000001", "0000001", "0000011", "0000001", "0000010", "0000001", "0000010", "0000000", "0000010", "0000001", "0000011", "0000001", "0000001", "0000010", "0000010", "0000011", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000010", "0000011", "0000000", "0000111", "0000010", "0000011", "0000010", "0000101", "0000011", "0001001", "0001000", "0001011", "0001011", "0000011", "0000110", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000011", "0000011", "0000001", "0000001", "0000011", "0000100", "0000100", "0000100", "0000000", "0000001", "0000010", "0000001", "0000001", "0000100", "0000001", "0000010", "0000010", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000010", "0000010", "0000100", "0000100", "0000001", "0000010", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000010", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000000", "0000010", "0000010", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000000", "0000010", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000000", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000010", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000010", "0000001", "0000001", "0000110", "0000010", "0000100", "0000010", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000010", "0000000", "0000001", "0000000", "0000010", "0000001", "0000011", "0000011", "0000101", "0000110", "0000010", "0000011", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0001000", "0001110", "0000111", "0001010", "0010011", "0000110", "0001101", "0001000", "0000001", "0000010", "0000100", "0000001", "0000011", "0000010", "0000011", "0000001", "0000010", "0000001", "0000101", "0000001", "0000010", "0000010", "0000011", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000100", "0000001", "0000011", "0000100", "0000000", "0001000", "0000011", "0000011", "0000010", "0000110", "0000011", "0001010", "0001001", "0001011", "0001010", "0000011", "0000110", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000010", "0000001", "0000010", "0000000", "0000101", "0000101", "0000010", "0000001", "0000101", "0000101", "0000110", "0000110", "0000100", "0001000", "0001111", "0000111", "0001001", "0010110", "0000111", "0001100", "0001001", "0000101", "0000100", "0001010", "0000011", "0000111", "0000100", "0001000", "0000010", "0000110", "0000101", "0001011", "0000010", "0000100", "0000111", "0000111", "0001010", "0000011", "0000101", "0000011", "0000110", "0000011", "0000100", "0000001", "0000010", "0000110", "0000010", "0000101", "0000010", "0000101", "0000010", "0000011", "0000100", "0000101", "0000101", "0000011", "0000100", "0001000", "0000010", "0000110", "0001001", "0000001", "0001011", "0000011", "0000100", "0000010", "0000110", "0000100", "0001001", "0001010", "0001101", "0001101", "0000100", "0001000", "0000111", "0000111", "0000011", "0000100", "0000011", "0000101", "0000101", "0000100", "0000011", "0000111", "0000111", "0000100", "0000110", "0000010", "0000010", "0000111", "0000100", "0000011", "0000111", "0000100", "0000011", "0001000", "0000101", "0000011", "0000110", "0010010", "0001100", "0000101", "0001100", "0000010", "0001110", "0010010", "0000110", "0000100", "0000111", "0000111", "0001010", "0001000", "0000101", "0001100", "0010110", "0001011", "0010000", "0010111", "0001000", "0001110", "0001001", "0000111", "0000100", "0001010", "0000011", "0000111", "0000101", "0001001", "0000011", "0000111", "0000111", "0001110", "0000011", "0000101", "0001000", "0001000", "0001011", "0000100", "0000111", "0000100", "0001001", "0000100", "0000101", "0000010", "0000010", "0001000", "0000011", "0001000", "0000011", "0000111", "0000011", "0000101", "0000110", "0000101", "0000110", "0000011", "0000100", "0001011", "0000011", "0001000", "0001011", "0000010", "0010001", "0000101", "0000110", "0000100", "0001000", "0000100", "0001101", "0001101", "0001100", "0001111", "0000100", "0000111", "0001101", "0001100", "0000100", "0000111", "0000101", "0001001", "0001000", "0000111", "0000101", "0001100", "0001101", "0000111", "0001010", "0000011", "0000100", "0001010", "0001000", "0000101", "0001100", "0000111", "0000110", "0001101", "0001000", "0000110", "0001011", "0010100", "0001110", "0000101", "0001110", "0000010", "0010000", "0010100", "0001000", "0000110", "0001011", "0001011", "0001111", "0001101", "0001000", "0000010", "0000101", "0000011", "0000011", "0000010", "0000010", "0000010", "0000001", "0001011", "0000010", "0000110", "0000010", "0000101", "0000011", "0000101", "0000010", "0000101", "0001010", "0001000", "0000010", "0000011", "0000111", "0000101", "0000111", "0000110", "0001010", "0000110", "0001101", "0000110", "0000111", "0000011", "0000100", "0001011", "0000101", "0001011", "0000100", "0001010", "0000100", "0000111", "0001000", "0000110", "0001000", "0000100", "0000101", "0001000", "0000010", "0000111", "0001001", "0000011", "0000110", "0000010", "0000010", "0000010", "0000001", "0000010", "0000010", "0000010", "0000001", "0000111", "0000001", "0000001", "0010010", "0010001", "0000110", "0001010", "0000111", "0001100", "0001011", "0001001", "0000110", "0010000", "0010010", "0001001", "0001110", "0000100", "0000110", "0010000", "0001010", "0001000", "0010010", "0001010", "0000111", "0010011", "0001100", "0001000", "0001111", "0011011", "0010100", "0000111", "0010100", "0000011", "0001111", "0010010", "0000111", "0000101", "0000100", "0000101", "0001001", "0000101", "0000011", "0000000", "0000001", "0000011", "0000001", "0000001", "0000010", "0000001", "0000001", "0000100", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000110", "0000001", "0000001", "0000010", "0000100", "0000010", "0000101", "0000010", "0000011", "0000001", "0000001", "0000100", "0000100", "0000100", "0000001", "0000100", "0000010", "0000011", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000010", "0000001", "0000001", "0000010", "0000111", "0000001", "0000010", "0001000", "0000111", "0000011", "0000101", "0000011", "0000101", "0000101", "0000100", "0000100", "0000111", "0001000", "0000101", "0000110", "0000010", "0000010", "0000110", "0000101", "0000011", "0000111", "0000100", "0000100", "0001000", "0000101", "0000011", "0001000", "0000101", "0000100", "0000001", "0000100", "0000010", "0000001", "0000010", "0000001", "0000011", "0000000", "0000010", "0000110", "0000001", "0000001", "0000010", "0000101", "0000011", "0000011", "0001001", "0000100", "0000110", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000110", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000011", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000010", "0000011", "0000000", "0000110", "0000010", "0000010", "0000010", "0000101", "0000100", "0001000", "0001001", "0001100", "0001111", "0000100", "0001000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000011", "0000001", "0000001", "0000110", "0000010", "0000010", "0000000", "0000010", "0000001", "0000001", "0000010", "0000001", "0000011", "0000001", "0000011", "0000110", "0000001", "0000100", "0010001", "0100000", "0010001", "0010101", "0101100", "0001110", "0011100", "0010001", "0000101", "0000100", "0001010", "0000011", "0000111", "0000100", "0001000", "0000011", "0000111", "0000101", "0001100", "0000100", "0000101", "0001011", "0001000", "0001010", "0000011", "0000101", "0000100", "0000110", "0000011", "0000100", "0000001", "0000010", "0000110", "0000101", "0000110", "0000010", "0000110", "0000010", "0000100", "0000100", "0000101", "0000110", "0000100", "0000101", "0001100", "0000011", "0001001", "0001100", "0000001", "0010011", "0000110", "0000111", "0000100", "0001011", "0000111", "0010011", "0010010", "0010111", "0010111", "0000111", "0001101", "0000100", "0000011", "0000001", "0000010", "0000100", "0000011", "0000010", "0000010", "0000100", "0000100", "0000100", "0000011", "0000011", "0000010", "0000001", "0000011", "0000010", "0000010", "0000011", "0000010", "0000101", "0000101", "0000011", "0000010", "0000111", "0001100", "0001001", "0000011", "0001000", "0000010", "0010000", "0010001", "0000111", "0000110", "0001100", "0001101", "0010001", "0001110", "0001010", "0000111", "0001101", "0001000", "0001001", "0001010", "0000101", "0000111", "0000101", "0001110", "0000110", "0010001", "0000101", "0001101", "0000111", "0001110", "0000101", "0001100", "0001110", "0010110", "0000101", "0001000", "0001101", "0001101", "0010010", "0000111", "0001100", "0001000", "0001111", "0001000", "0001001", "0000100", "0000101", "0001110", "0000111", "0001111", "0000110", "0001101", "0000110", "0001001", "0001010", "0001010", "0001011", "0000110", "0001000", "0010010", "0000101", "0001110", "0010011", "0000100", "0011001", "0000111", "0001001", "0000110", "0001011", "0000111", "0010001", "0010010", "0010000", "0010010", "0000101", "0001010", "0011010", "0010111", "0001001", "0001110", "0001001", "0010001", "0010000", "0001100", "0001001", "0010111", "0011010", "0001101", "0010011", "0000101", "0001000", "0010110", "0001110", "0001011", "0011000", "0001110", "0001010", "0011001", "0010001", "0001100", "0010101", "0100110", "0011100", "0001011", "0011100", "0000100", "0011000", "0011111", "0001100", "0001001", "0001010", "0001011", "0010001", "0001100", "0001001", "0000100", "0000111", "0000110", "0000100", "0001100", "0000110", "0000111", "0000101", "0001101", "0000100", "0001001", "0000011", "0000111", "0000100", "0001000", "0000100", "0000110", "0001100", "0001101", "0000100", "0000101", "0001011", "0001000", "0001011", "0000111", "0001100", "0001000", "0001111", "0000111", "0001000", "0000100", "0000100", "0001101", "0000111", "0001101", "0000101", "0001100", "0000101", "0001000", "0001010", "0000110", "0001000", "0000100", "0000101", "0001001", "0000011", "0000111", "0001001", "0000100", "0001100", "0000100", "0000101", "0000011", "0000110", "0000101", "0001100", "0001010", "0001101", "0001111", "0000100", "0001000", "0001011", "0001001", "0000100", "0000111", "0001000", "0000111", "0000111", "0000110", "0000111", "0001010", "0001011", "0000110", "0001001", "0000101", "0000011", "0001010", "0000110", "0000101", "0001011", "0000110", "0001010", "0001011", "0000111", "0000101", "0001101", "0001010", "0001000", "0000011", "0000111", "0000100", "0000101", "0000110", "0000010", "0000110", "0000010", "0000110", "0001011", "0000011", "0000111", "0010010", "0100001", "0010010", "0011000", "0101101", "0001110", "0011100", "0010001", "0001001", "0001011", "0011010", "0001000", "0010011", "0001011", "0010110", "0000111", "0010011", "0001000", "0100001", "0000111", "0001100", "0010010", "0010100", "0011011", "0000101", "0001000", "0000101", "0001011", "0000101", "0000110", "0000011", "0000011", "0001010", "0000110", "0001001", "0000011", "0001001", "0000100", "0000110", "0000110", "0000111", "0000111", "0000100", "0000101", "0001100", "0000100", "0001001", "0001101", "0000010", "0010010", "0000101", "0000110", "0000100", "0001011", "0000111", "0010001", "0010001", "0010110", "0010111", "0000111", "0001100", "0001010", "0001001", "0000011", "0000101", "0000110", "0000111", "0000110", "0000101", "0000110", "0001001", "0001010", "0000101", "0000111", "0000100", "0000011", "0001000", "0000110", "0000101", "0001010", "0000110", "0001000", "0001100", "0000111", "0000101", "0001100", "0010111", "0010001", "0000110", "0010000", "0000011", "0010111", "0011011", "0001010", "0001000", "0001110", "0010001", "0011000", "0010001", "0001101", "0000100", "0001000", "0000101", "0000101", "0000101", "0000011", "0000011", "0000010", "0010010", "0000011", "0001000", "0000011", "0000110", "0000011", "0000110", "0000011", "0000101", "0010000", "0001000", "0000011", "0000101", "0001011", "0000110", "0000110", "0001010", "0010001", "0001011", "0010101", "0001010", "0001011", "0000101", "0000111", "0010010", "0001001", "0010010", "0000111", "0010001", "0000111", "0001011", "0001100", "0001110", "0001111", "0001000", "0001011", "0011011", "0000111", "0010100", "0011100", "0000101", "0101000", "0001100", "0001111", "0001001", "0010110", "0001101", "0100010", "0100011", "0100101", "0100110", "0001100", "0010111", "0011011", "0010111", "0001001", "0001111", "0001010", "0010001", "0010000", "0001110", "0001010", "0011000", "0011010", "0001101", "0010101", "0000111", "0001000", "0010111", "0001111", "0001011", "0011010", "0001111", "0001100", "0011001", "0010001", "0001100", "0010111", "0100000", "0010110", "0001000", "0010111", "0000101", "0010001", "0010101", "0001001", "0001000", "0000110", "0000111", "0001110", "0001000", "0010001", "0000000", "0000010", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0010110", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0010110", "0000001", "0000010", "0000011", "0001110", "0000010", "0000001", "0001100", "0010110", "0001101", "0011011", "0001101", "0001111", "0000110", "0001000", "0010111", "0001100", "0011000", "0001000", "0010101", "0001001", "0001110", "0010001", "0001100", "0001111", "0001000", "0001010", "0010001", "0000101", "0001101", "0010010", "0000111", "0010010", "0000101", "0000110", "0000100", "0000111", "0000101", "0001011", "0001011", "0001001", "0001100", "0000011", "0000110", "0000011", "0000010", "0000001", "0000010", "0001110", "0000010", "0000010", "0000010", "0001000", "0000011", "0000010", "0000011", "0000010", "0001001", "0000001", "0000010", "0000010", "0000010", "0000011", "0000011", "0001111", "0001000", "0000011", "0000001", "0001110", "0000110", "0000010", "0000001", "0000011", "0000111", "0000001", "0000001", "0000001", "0001000", "0000001", "0000010", "0001101", "0000001", "0000100", "0000000", "0000010", "0000010", "0000000", "0000000", "0000010", "0000000", "0000000", "0000011", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000011", "0000001", "0000001", "0000011", "0010100", "0000011", "0000001", "0000011", "0000011", "0000010", "0000100", "0000011", "0000011", "0000010", "0000001", "0000100", "0001101", "0000100", "0000001", "0000011", "0000001", "0000011", "0000011", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000111", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000001", "0000010", "0001010", "0000010", "0000001", "0000010", "0000001", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0001010", "0001001", "0000011", "0000001", "0010001", "0000110", "0000001", "0000000", "0000010", "0000010", "0000000", "0000001", "0000000", "0001010", "0000000", "0000010", "0010000", "0000000", "0000101", "0000000", "0000011", "0000010", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000011", "0010101", "0000110", "0000001", "0000010", "0000001", "0000000", "0000001", "0000010", "0000010", "0000001", "0000001", "0000010", "0001110", "0000001", "0000000", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000111", "0000011", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0001100", "0000011", "0000001", "0000010", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0001111", "0001010", "0000011", "0000001", "0010010", "0000111", "0000001", "0000000", "0000010", "0000011", "0000001", "0000001", "0000000", "0001011", "0000000", "0000010", "0011011", "0000000", "0000111", "0000000", "0000100", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000011", "0000010", "0000001", "0000000", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000100", "0010011", "0000101", "0000001", "0000010", "0000001", "0000000", "0000001", "0000100", "0000011", "0000010", "0000001", "0000010", "0001100", "0000001", "0000000", "0000001", "0000001", "0000010", "0000011", "0000001", "0000001", "0000000", "0000001", "0000011", "0000001", "0000001", "0000001", "0000000", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000111", "0000100", "0000100", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000101", "0001011", "0000100", "0000001", "0000010", "0000001", "0000110", "0000001", "0000001", "0000001", "0000010", "0000001", "0000100", "0001111", "0001001", "0000011", "0000001", "0010001", "0000110", "0000001", "0000000", "0000011", "0000011", "0000001", "0000001", "0000000", "0001011", "0000001", "0000010", "0010110", "0000000", "0001100", "0000000", "0000111", "0000011", "0000001", "0000001", "0000010", "0000001", "0000001", "0000110", "0000100", "0000100", "0000011", "0000001", "0000000", "0000001", "0000010", "0000001", "0000110", "0000001", "0000001", "0000100", "0011011", "0000101", "0000001", "0000101", "0000110", "0000100", "0001000", "0000110", "0000101", "0000011", "0000010", "0000111", "0010001", "0000111", "0000010", "0000110", "0000010", "0000101", "0000111", "0000100", "0000101", "0000011", "0000100", "0001011", "0000011", "0001000", "0001010", "0000010", "0010000", "0000101", "0000110", "0000100", "0000101", "0000100", "0001001", "0001001", "0010100", "0010111", "0001000", "0001110", "0000001", "0000001", "0000001", "0000001", "0000100", "0000010", "0000001", "0000111", "0010000", "0000100", "0000001", "0000010", "0000001", "0000111", "0000001", "0000001", "0000010", "0000010", "0000001", "0000101", "0010010", "0001100", "0000100", "0000010", "0010111", "0001000", "0000001", "0000000", "0000011", "0000100", "0000001", "0000001", "0000000", "0001110", "0000001", "0000010", "0010111", "0000001", "0011000", "0000111", "0001110", "0000111", "0001001", "0001111", "0000101", "0001001", "0000110", "0100000", "0000101", "0000101", "0000011", "0000010", "0000001", "0000011", "0000011", "0000010", "0011110", "0000011", "0000010", "0000110", "0100110", "0001010", "0000100", "0010001", "0011110", "0010011", "0100110", "0010011", "0010101", "0001010", "0001011", "0100001", "0011101", "0100010", "0001101", "0100000", "0001101", "0010110", "0011001", "0010111", "0011011", "0001111", "0010011", "0100100", "0001010", "0011100", "0100111", "0001001", "0101111", "0001110", "0010001", "0001011", "0011001", "0001111", "0101001", "0101010", "0100101", "0101000", "0001111", "0011010", "0000101", "0000101", "0000010", "0000011", "0010100", "0000100", "0000011", "0000111", "0011100", "0001000", "0000101", "0000011", "0000100", "0001110", "0000010", "0000100", "0000100", "0000011", "0000101", "0000111", "0100010", "0010101", "0001001", "0000011", "0101010", "0010011", "0000110", "0000010", "0001000", "0001011", "0001000", "0001001", "0000100", "0010110", "0000100", "0000101", "0101010", "0000101", "0011010", "0101011", "1010100", "0101010", "0111000", "1011011", "0100000", "0111010", "0100101", "0011110", "0010100", "0101101", "0001111", "0100000", "0010011", "0100100", "0001100", "0011110", "0011100", "0111010", "0001101", "0010111", "0111110", "0100111", "0110000", "0010001", "0011110", "0010011", "0100101", "0010100", "0010011", "0001001", "0001011", "0100001", "0101100", "0011111", "0001101", "0100000", "0001101", "0010110", "0010111", "0010011", "0010111", "0001100", "0010000", "0100010", "0001010", "0011010", "0100011", "0001001", "0101010", "0001100", "0001111", "0001001", "0011000", "0010001", "0101000", "0100111", "0011100", "0011101", "0001110", "0010110", "1000011", "0111100", "0010111", "0100110", "0010101", "0101111", "0101001", "0100010", "0101011", "0111110", "1000001", "0100001", "0110100", "0010000", "0010101", "0111011", "0101000", "0011101", "1000010", "0101000", "0101100", "1000111", "0101110", "0100000", "1010101", "1101101", "1010001", "0011110", "1010000", "0001011", "1001010", "1011011", "0100011", "0101101", "0101000", "0101100", "1011000", "0110010", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0001010", "0000101", "0000101", "0000000", "0001010", "0000101", "0001010", "0000101", "0011001", "0000000", "0001010", "0001010", "0001010", "0000101", "0000000", "0000101", "0001010", "0000101", "0000000", "0011110", "0000101", "0100011", "0001010", "0001111", "0010100", "0000000", "0000000", "0000000", "0000000", "0000101", "0000000", "0000000", "0000000", "0001010", "0000000", "0000101", "0000101", "0011001", "0001010", "0001010", "0000101", "0000101", "0000101", "0000000", "0000000", "0000000", "0000000", "0000000", "0011001", "0001111", "0001010", "0010100", "0011110", "0001111", "0000101", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000101", "0001010", "0000101", "0000101", "0000101", "0000101", "0000101", "0000101", "0000101", "0000101", "0001111", "0000101", "0000101", "0011001", "0000000", "0000101", "0000000", "0011001", "0011001", "0001111", "0001010", "0000000", "0001111", "0010100", "0000000", "0000000", "0000000", "0001101", "0000110", "0001011", "0010010", "0001010", "0010010", "0011000", "0011110", "0011111", "0010100", "0010101", "0010101", "0011001", "0010011", "0011011", "0010001", "0110010", "0001110", "0101100", "0010011", "0110010", "0100110", "0011011", "0100110", "0110100", "0100010", "0001101", "0101101", "0010000", "0110001", "0100111", "0101000", "0110000", "0111110", "0101111", "0100010", "0100001", "0110101", "0100100", "0010001", "0010111", "0100000", "0001010", "0001110", "0010000", "0100011", "0011111", "0011100", "0010111", "0011001", "0011101", "0011010", "0010000", "0001000", "0010101", "0000110", "0100100", "0011001", "0001111", "0100010", "0100001", "0101110", "0001010", "0010110", "0001010", "0001000", "0001101", "0010001", "0010101", "0011000", "0001111", "0001101", "0001001", "0010010", "0010010", "0001101", "0001110", "0010011", "0001010", "0001011", "0001011", "0010110", "0010011", "0101100", "0010010", "0010010", "0100100", "0001100", "0011100", "0001101", "0111010", "0011010", "0111110", "0011000", "0001001", "0011000", "0011010", "0010100", "0011101", "0011011", "0001111", "0000110", "0001100", "0010110", "0001110", "0010101", "0011010", "0100000", "0100001", "0010110", "0010111", "0010111", "0010110", "0010100", "0011011", "0010001", "0110101", "0001111", "0110000", "0010000", "0110010", "0100111", "0011011", "0101010", "0110110", "0100110", "0001100", "0101010", "0001101", "0101110", "0110001", "0110000", "0111011", "0101001", "0011110", "0010110", "0110000", "1001010", "0110111", "0010100", "0011011", "0100001", "0001011", "0001110", "0010000", "0011001", "0010111", "0001101", "0010011", "0010101", "0011000", "0010101", "0001111", "0000111", "0010011", "0000101", "0100010", "0011001", "0001111", "0100010", "0100010", "0100010", "0001000", "0010010", "0001000", "0000110", "0001101", "0010001", "0010111", "0100010", "0010001", "0010010", "0001000", "0010000", "0010000", "0001100", "0001101", "0010010", "0001000", "0001001", "0001001", "0010011", "0010000", "0101100", "0010000", "0010000", "0100000", "0001010", "0011100", "0001101", "1000100", "0011101", "0111001", "0010100", "0000111", "0010110", "0011000", "0010001", "0011000", "0010101", "0001111", "0001000", "0001100", "0100010", "0010010", "0100011", "0101110", "0110110", "0111000", "0100101", "0100111", "0100001", "0101111", "0100001", "0101111", "0011110", "0100111", "0010111", "1001110", "0100011", "1010111", "1000011", "0101111", "1001100", "1100100", "1000011", "0011000", "1001110", "0010111", "1010110", "1000010", "1000011", "1010000", "1110100", "1010110", "1000010", "0111000", "1001110", "0111101", "0101011", "0110111", "1000010", "0010000", "0010100", "0011000", "0111100", "0110110", "0010110", "0101001", "0101110", "0110100", "0101101", "0011111", "0001111", "0100011", "0001011", "0111111", "0101001", "0011010", "0110111", "0110110", "0110100", "0010011", "0100001", "0001111", "0001011", "0001110", "0010001", "0010101", "0101111", "0010110", "0011010", "0010000", "0100010", "0100001", "0011001", "0011001", "0100011", "0001111", "0010011", "0010100", "0101001", "0100010", "0110110", "0100000", "0011111", "0101001", "0010100", "0111001", "0011000", "1000001", "0110011", "0101111", "0101100", "0001100", "0101100", "0101011", "0011101", "0101100", "0100110", "0101100", "0010101", "0011111", "1000110", "0100100", "1000111", "0010001", "0010101", "0010100", "0001110", "0001111", "0001101", "0111001", "0001101", "0010011", "0001011", "0010001", "0001001", "0011101", "0101011", "0100001", "0011010", "0010010", "0011101", "0100111", "0011010", "0011101", "0100110", "0001100", "0101011", "0100111", "0100110", "0110001", "0101001", "0100000", "0010111", "0101010", "0110110", "0101110", "0011001", "0100001", "0101010", "0011101", "0100101", "0101000", "1001011", "1000000", "0011010", "0110100", "0111000", "0111110", "0110111", "0101000", "0010001", "0101100", "0001101", "1100001", "1000001", "0101001", "1010111", "1010111", "1010010", "0010101", "0110010", "0010110", "0010001", "0100010", "0110110", "0111110", "1011001", "0100101", "0110010", "0010011", "0101000", "0101001", "0011101", "0100000", "0101100", "0010001", "0010111", "0011001", "0110001", "0101011", "0111110", "0101000", "0101001", "0101011", "0011100", "1001000", "0100000", "1010111", "1010001", "0110101", "0110011", "0010101", "1000110", "1001010", "0110100", "1001000", "1000000", "0001001", "0000100", "0000111", "0001101", "0000111", "0001110", "0010010", "0010110", "0011000", "0001111", "0010000", "0001110", "0101110", "0001110", "0010100", "0001100", "0010001", "0001010", "0100010", "0100000", "0100100", "0011100", "0010011", "0011111", "0101011", "0011011", "0010110", "0100000", "0001010", "0100100", "0011110", "0011111", "0100100", "0100111", "0011110", "0010101", "0011010", "0100010", "0011100", "0001010", "0001110", "0010001", "0001001", "0001011", "0001110", "0111000", "0110011", "0010101", "0100100", "0101001", "0101110", "0101001", "0011110", "0001110", "0100000", "0001010", "0111110", "0101001", "0011010", "0110110", "0110101", "0110011", "0010001", "0011111", "0001110", "0001010", "0010010", "0011001", "0011100", "0011110", "0001101", "0010000", "0000101", "0001100", "0001011", "0001001", "0001001", "0001100", "0000101", "0010001", "0000111", "0001111", "0001100", "0010101", "0001011", "0001100", "0100000", "0000111", "0010100", "0001001", "0011000", "0010010", "0010110", "0101001", "0000101", "0001111", "0010000", "0001100", "0010010", "0010000", "0010000", "0001000", "0001100", "0010110", "0001100", "0010111", "0001110", "0010010", "0010001", "0001100", "0001101", "0001010", "0100000", "0001011", "0010001", "0001001", "0010001", "0000111", "0011000", "0011000", "0011100", "0010110", "0001111", "0011001", "0011111", "0010110", "0010000", "0011101", "0001001", "0100000", "0011111", "0011111", "0100111", "0101011", "0100010", "0011001", "0011100", "0100101", "0011111", "0010010", "0010110", "0011100", "0010010", "0011000", "0011010", "0101010", "0100011", "0001110", "0011011", "0011110", "0100010", "0011110", "0010101", "0001001", "0011000", "0001000", "0111011", "0100111", "0011000", "0111101", "0111100", "0111001", "0001011", "0101000", "0010011", "0001101", "0011000", "0100101", "0101001", "1000110", "0011110", "0100110", "0010001", "0100010", "0100100", "0011011", "0011101", "0100101", "0001110", "0001101", "0010110", "0101011", "0100011", "0110011", "0100011", "0100100", "0011000", "0010111", "0111011", "0011011", "0111111", "0111010", "0101100", "0011101", "0001110", "0101110", "0110010", "0011110", "0101110", "0101000", "0100010", "0010000", "0011001", "1000011", "0100010", "1000100", "0000110", "0000111", "0001000", "0000101", "0000110", "0000110", "0001000", "0000100", "0001010", "0000100", "0001011", "0000100", "0001011", "0000110", "0001100", "0001010", "0000110", "0001001", "0001111", "0001001", "0000101", "0001101", "0000100", "0001110", "0001100", "0001101", "0001111", "0010110", "0010001", "0001001", "0010101", "0011010", "0010101", "0001101", "0010001", "0010101", "0000110", "0001000", "0001001", "0001011", "0001010", "0000100", "0000111", "0001000", "0001001", "0000111", "0000101", "0000011", "0000110", "0000010", "0001101", "0001000", "0000101", "0001110", "0001110", "0001101", "0000011", "0001011", "0000101", "0000100", "0001011", "0001100", "0001111", "0011111", "0001101", "0010010", "0001011", "0010110", "0010111", "0010001", "0010010", "0011001", "0001010", "0000100", "0001110", "0011110", "0011000", "0100100", "0011000", "0010101", "0001100", "0001111", "0101000", "0010001", "0110110", "0101101", "0100011", "0001000", "0001101", "0101010", "0101011", "0101000", "0110110", "0110001", "0010000", "0000111", "0001011", "0011011", "0001100", "0010111", "0000101", "0000110", "0000110", "0000100", "0000100", "0000100", "0000110", "0000100", "0001000", "0000011", "0001011", "0000011", "0001001", "0000101", "0001010", "0000111", "0000101", "0001000", "0001001", "0001000", "0000100", "0001001", "0000011", "0001011", "0001001", "0001001", "0001011", "0010011", "0001111", "0001000", "0001011", "0001101", "0001010", "0000100", "0000111", "0001000", "0000011", "0000100", "0000101", "0000111", "0000111", "0000011", "0000101", "0000110", "0000111", "0000110", "0000100", "0000010", "0000101", "0000001", "0001010", "0000110", "0000100", "0001010", "0001000", "0001000", "0000010", "0000110", "0000010", "0000010", "0001000", "0000110", "0000111", "0001010", "0000100", "0000101", "0000110", "0001011", "0001011", "0001001", "0001001", "0001101", "0000101", "0000011", "0000111", "0001111", "0001100", "0010010", "0001100", "0001100", "0000110", "0000111", "0010101", "0001001", "0011010", "0010110", "0010010", "0000110", "0000111", "0010111", "0010111", "0010011", "0011000", "0010100", "0000111", "0000100", "0000101", "0001101", "0001010", "0010010", "0000100", "0000100", "0000101", "0000011", "0000011", "0000011", "0000111", "0000011", "0001000", "0000010", "0001000", "0000011", "0000110", "0000101", "0000111", "0000111", "0000100", "0000110", "0001000", "0000110", "0000100", "0000110", "0000010", "0000111", "0000110", "0000111", "0001001", "0010000", "0001110", "0000111", "0001011", "0001010", "0001010", "0000101", "0000111", "0001001", "0000011", "0000100", "0000100", "0001001", "0001000", "0000100", "0000110", "0000111", "0001000", "0000111", "0000101", "0000010", "0000101", "0000010", "0001001", "0001000", "0000101", "0001001", "0001010", "0001010", "0000011", "0000101", "0000011", "0000010", "0001000", "0000100", "0000101", "0001001", "0000101", "0000110", "0000001", "0000011", "0000011", "0000010", "0000010", "0000100", "0000010", "0000011", "0000010", "0000011", "0000100", "0000111", "0000011", "0000011", "0000110", "0000010", "0000101", "0000010", "0001100", "0000111", "0001001", "0000111", "0000010", "0001001", "0001001", "0000110", "0001110", "0001010", "0000100", "0000001", "0000001", "0000010", "0000011", "0000010", "0000100", "0000100", "0000100", "0000011", "0000011", "0000011", "0000010", "0000011", "0000111", "0000010", "0000111", "0000100", "0000110", "0000001", "0000110", "0000111", "0000011", "0000101", "0000111", "0000100", "0000011", "0000110", "0000010", "0000111", "0000110", "0000110", "0000111", "0001110", "0001101", "0000101", "0001010", "0001000", "0000111", "0000100", "0000110", "0000110", "0000010", "0000010", "0000011", "0000010", "0000010", "0000010", "0000010", "0000010", "0000010", "0000011", "0000001", "0000001", "0000010", "0000000", "0000101", "0000101", "0000010", "0000100", "0000110", "0000101", "0000001", "0000100", "0000011", "0000010", "0001000", "0000110", "0000110", "0000111", "0000101", "0000101", "0000001", "0000011", "0000011", "0000010", "0000010", "0000100", "0000001", "0000001", "0000010", "0000011", "0000110", "0000110", "0000011", "0000011", "0000100", "0000010", "0000101", "0000010", "0001010", "0000011", "0001000", "0000010", "0000001", "0000010", "0000010", "0000010", "0000010", "0000010", "0000100", "0000010", "0000010", "0000100", "0000100", "0000011", "0000011", "0000011", "0000011", "0000010", "0000010", "0000011", "0000101", "0000011", "0000111", "0000010", "0001000", "0000100", "0000100", "0000100", "0000100", "0000111", "0000010", "0000100", "0000101", "0000011", "0000100", "0000101", "0000010", "0000110", "0000101", "0000110", "0001000", "0001111", "0001101", "0000101", "0001001", "0001001", "0000111", "0000100", "0000110", "0000110", "0000100", "0000101", "0000110", "0000110", "0000101", "0000010", "0000101", "0000100", "0000101", "0000101", "0000011", "0000001", "0000011", "0000001", "0000100", "0000110", "0000010", "0000011", "0000010", "0000011", "0000010", "0000001", "0000001", "0000001", "0000111", "0000001", "0000001", "0000011", "0000010", "0000001", "0000101", "0001001", "0001010", "0000111", "0000111", "0001010", "0000100", "0000010", "0000101", "0001011", "0001011", "0001110", "0001001", "0001001", "0000110", "0000110", "0010000", "0000111", "0010001", "0001111", "0001100", "0000100", "0000011", "0001001", "0001010", "0000110", "0000111", "0000110", "0001010", "0000101", "0000111", "0001111", "0001001", "0010001", "0000111", "0001001", "0001001", "0000101", "0000110", "0000110", "0001011", "0000110", "0001011", "0000101", "0001000", "0000101", "0001101", "0001000", "0001110", "0001100", "0000111", "0001100", "0001111", "0001010", "0000110", "0001001", "0000010", "0001001", "0000110", "0000110", "0000111", "0001100", "0001101", "0000011", "0001000", "0000110", "0000101", "0000010", "0000101", "0000101", "0000100", "0000101", "0000101", "0001101", "0001100", "0000101", "0001001", "0001010", "0001011", "0001010", "0000111", "0000011", "0000111", "0000010", "0010000", "0001011", "0000111", "0001100", "0001110", "0001100", "0000100", "0000111", "0000011", "0000010", "0001000", "0000100", "0000101", "0000101", "0000010", "0000011", "0000110", "0001100", "0001011", "0001001", "0001001", "0001100", "0000101", "0000100", "0000111", "0001101", "0001100", "0010001", "0001011", "0001011", "0001000", "0001000", "0010011", "0001001", "0010111", "0010100", "0001110", "0001010", "0000101", "0010001", "0010010", "0001011", "0010011", "0010000", "0001011", "0000101", "0001000", "0010100", "0001011", "0010100", "0000111", "0000111", "0001000", "0000110", "0000110", "0000100", "0001011", "0000101", "0001010", "0000100", "0000110", "0000100", "0001011", "0001000", "0001100", "0001010", "0000110", "0001010", "0001101", "0001001", "0000110", "0010001", "0000101", "0010010", "0010011", "0010011", "0010110", "0011001", "0010110", "0001111", "0010001", "0010100", "0010000", "0000111", "0001001", "0001010", "0000010", "0000011", "0000011", "0001110", "0001101", "0000101", "0001010", "0001010", "0001101", "0001011", "0000111", "0000011", "0001001", "0000011", "0010010", "0001100", "0000111", "0010001", "0010000", "0001111", "0000100", "0001001", "0000101", "0000011", "0001010", "0001010", "0001010", "0010001", "0001000", "0001010", "0000001", "0000011", "0000011", "0000010", "0000010", "0000100", "0000010", "0000100", "0000010", "0000100", "0000100", "0000110", "0000011", "0000100", "0001001", "0000010", "0000101", "0000011", "0001100", "0001010", "0001010", "0001010", "0000100", "0001101", "0001100", "0001101", "0010011", "0010001", "0000100", "0000010", "0000010", "0001010", "0000101", "0001010", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000111", "0000001", "0000011", "0000010", "0000001", "0000010", "0000010", "0000011", "0000001", "0000010", "0000010", "0000001", "0000011", "0000011", "0000001", "0000011", "0000101", "0000101", "0000110", "0010100", "0001111", "0000111", "0010000", "0010011", "0010001", "0001100", "0001111", "0010011", "0000001", "0000001", "0000001", "0000100", "0000100", "0000010", "0000011", "0000011", "0000011", "0000100", "0000010", "0000001", "0000011", "0000001", "0000111", "0000110", "0000011", "0001011", "0001011", "0001010", "0000001", "0001010", "0000100", "0000011", "0001001", "0001011", "0001101", "0010100", "0001000", "0001100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000010", "0000001", "0000001", "0000010", "0000011", "0000001", "0000010", "0000100", "0000001", "0000001", "0000001", "0000110", "0000001", "0000110", "0000011", "0000001", "0000001", "0000001", "0000010", "0000011", "0000011", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000110", "0000010", "0000111", "0000001", "0000100", "0000010", "0000010", "0000101", "0000010", "0000010", "0000001", "0000001", "0000010", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0001011", "0001100", "0000001", "0000111", "0000011", "0000010", "0000010", "0000011", "0000011", "0000011", "0000100", "0000100", "0001000", "0000110", "0000011", "0000110", "0000110", "0000110", "0000110", "0000100", "0000010", "0000101", "0000001", "0000101", "0000100", "0000010", "0000011", "0000011", "0000011", "0000010", "0000010", "0000001", "0000001", "0000111", "0000011", "0000100", "0001010", "0000011", "0000101", "0000001", "0000010", "0000011", "0000010", "0000010", "0000011", "0000001", "0000011", "0000001", "0000011", "0000011", "0000101", "0000010", "0000011", "0000101", "0000010", "0000100", "0000010", "0000110", "0000010", "0000110", "0000110", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000110", "0000111", "0000111", "0000101", "0000101", "0000100", "0001110", "0000100", "0001001", "0000100", "0000101", "0000011", "0001001", "0001010", "0001010", "0001000", "0000110", "0001001", "0001100", "0001000", "0000111", "0000111", "0000010", "0001000", "0000011", "0000100", "0000101", "0001100", "0001100", "0000010", "0000111", "0000010", "0000010", "0000001", "0000010", "0000001", "0000100", "0000110", "0000110", "0010001", "0001111", "0000110", "0001100", "0001101", "0001111", "0001101", "0001001", "0000100", "0001010", "0000011", "0010100", "0001101", "0001001", "0001111", "0001111", "0001110", "0000101", "0000101", "0000010", "0000010", "0000111", "0000011", "0000100", "0000011", "0000010", "0000010", "0000101", "0001011", "0001100", "0001000", "0001001", "0001100", "0000100", "0000110", "0000111", "0001110", "0001100", "0010001", "0001011", "0001011", "0001010", "0000111", "0010100", "0001001", "0010001", "0001111", "0001011", "0001100", "0000010", "0001000", "0001000", "0000011", "0000100", "0000100", "0001001", "0000100", "0000110", "0001011", "0000110", "0001011", "0000100", "0000101", "0000101", "0000011", "0000011", "0000011", "0001000", "0000011", "0001000", "0000010", "0000101", "0000010", "0000110", "0000110", "0000111", "0000110", "0000100", "0000111", "0001001", "0000110", "0000101", "0001010", "0000011", "0001011", "0001100", "0001011", "0001110", "0010010", "0010000", "0001000", "0001011", "0001010", "0001000", "0000011", "0000100", "0000101", "0000011", "0000100", "0000101", "0001011", "0001001", "0000011", "0000111", "0001000", "0001001", "0001000", "0000110", "0000010", "0000110", "0000010", "0001100", "0001001", "0000110", "0010000", "0001111", "0001110", "0000011", "0001101", "0000110", "0000100", "0001010", "0001100", "0001110", "0010101", "0000111", "0001100", "0000100", "0001001", "0001001", "0000111", "0000111", "0001010", "0000100", "0000011", "0000110", "0001011", "0001010", "0001110", "0001001", "0001001", "0000110", "0000110", "0010000", "0000110", "0010100", "0010001", "0001100", "0000111", "0000110", "0010001", "0010010", "0001110", "0010101", "0010000", "0001010", "0000101", "0000111", "0010011", "0001011", "0010100", "0000100", "0000100", "0000100", "0000011", "0000011", "0000010", "0000110", "0000010", "0000101", "0000010", "0000011", "0000010", "0000110", "0000101", "0000110", "0000101", "0000011", "0000110", "0000111", "0000101", "0000011", "0000110", "0000010", "0000110", "0000110", "0000110", "0000110", "0001011", "0001001", "0000110", "0001100", "0001111", "0001100", "0001000", "0001011", "0001101", "0000001", "0000010", "0000010", "0001000", "0000111", "0000011", "0000101", "0000110", "0000111", "0000110", "0000100", "0000010", "0000101", "0000001", "0001011", "0001000", "0000101", "0001100", "0001100", "0001011", "0000010", "0000111", "0000011", "0000010", "0000101", "0000111", "0001000", "0010000", "0000111", "0001001", "0000011", "0000101", "0000101", "0000100", "0000100", "0000110", "0000010", "0000010", "0000011", "0000111", "0000110", "0001000", "0000101", "0000101", "0000100", "0000100", "0001001", "0000100", "0001100", "0001100", "0001000", "0000110", "0000100", "0001100", "0001100", "0001010", "0001111", "0001101", "0000110", "0000011", "0000101", "0001110", "0000111", "0001101", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000010", "0000011", "0000010", "0000001", "0000100", "0000001", "0000101", "0000110", "0000110", "0001000", "0001001", "0000110", "0000100", "0000101", "0000111", "0000110", "0000100", "0000100", "0000101", "0000000", "0000000", "0000000", "0000011", "0000010", "0000001", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000010", "0000000", "0000101", "0000011", "0000010", "0000110", "0000111", "0000111", "0000001", "0000110", "0000011", "0000010", "0000100", "0000111", "0001000", "0001110", "0000101", "0001000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000100", "0000011", "0000010", "0000010", "0000010", "0000110", "0000110", "0000111", "0001010", "0001000", "0000010", "0000001", "0000001", "0000111", "0000011", "0000111", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000100", "0000011", "0000011", "0000110", "0000111", "0000110", "0000100", "0000101", "0000111", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000010", "0000010", "0000010", "0000000", "0000010", "0000001", "0000001", "0000010", "0000011", "0000100", "0001000", "0000011", "0000101", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000010", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000010", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000000", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000011", "0000010", "0000010", "0000010", "0000011", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000010", "0000100", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000010", "0000010", "0001001", "0000100", "0001001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000010", "0000010", "0000011", "0000110", "0000100", "0000011", "0000110", "0001001", "0000111", "0000101", "0000110", "0000111", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000010", "0000001", "0000001", "0000011", "0000011", "0000011", "0000000", "0000011", "0000001", "0000001", "0000010", "0000100", "0000100", "0001010", "0000100", "0000101", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000010", "0000010", "0000111", "0000011", "0000101", "0001101", "0000111", "0001101", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000011", "0000001", "0000010", "0000001", "0000001", "0000001", "0000011", "0000010", "0000011", "0000011", "0000010", "0000011", "0000100", "0000011", "0000001", "0000110", "0000010", "0000110", "0000111", "0000110", "0001000", "0001000", "0000110", "0000100", "0000101", "0000111", "0000110", "0000100", "0000101", "0000110", "0000000", "0000000", "0000000", "0000011", "0000011", "0000001", "0000010", "0000011", "0000011", "0000010", "0000010", "0000001", "0000010", "0000001", "0000110", "0000100", "0000011", "0001001", "0001000", "0001000", "0000001", "0000111", "0000011", "0000010", "0000100", "0000111", "0001000", "0001100", "0000101", "0000111", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000101", "0000101", "0000011", "0000010", "0000010", "0000111", "0001000", "0001000", "0001100", "0001010", "0001011", "0000101", "0000111", "0010110", "0001010", "0010110", "0000100", "0000100", "0000100", "0000011", "0000011", "0000010", "0000111", "0000010", "0000101", "0000010", "0000011", "0000010", "0000101", "0000101", "0000110", "0000101", "0000011", "0000101", "0000111", "0000100", "0000100", "0000101", "0000010", "0000110", "0000110", "0000110", "0001000", "0001110", "0001011", "0000111", "0001110", "0010000", "0001101", "0001000", "0001010", "0001101", "0000010", "0000010", "0000010", "0001001", "0001000", "0000011", "0000111", "0000111", "0001000", "0000111", "0000101", "0000010", "0000101", "0000010", "0001100", "0001000", "0000101", "0001011", "0001011", "0001011", "0000011", "0000111", "0000011", "0000010", "0000111", "0001000", "0001001", "0010101", "0001000", "0001100", "0000011", "0000110", "0000111", "0000101", "0000101", "0000111", "0000011", "0000011", "0000100", "0001000", "0000111", "0001001", "0000110", "0000110", "0000101", "0000100", "0001011", "0000101", "0001110", "0001101", "0001001", "0000111", "0000100", "0001100", "0001110", "0001100", "0010000", "0001101", "0000110", "0000011", "0000101", "0000111", "0000101", "0000111", "0000101", "0000110", "0000110", "0000100", "0000100", "0000011", "0001000", "0000011", "0001001", "0000011", "0000101", "0000011", "0001000", "0000110", "0001001", "0001000", "0000101", "0001000", "0001010", "0000111", "0000101", "0001011", "0000011", "0001101", "0001100", "0001011", "0001101", "0010001", "0010000", "0000111", "0001001", "0001000", "0000110", "0000010", "0000011", "0000011", "0000100", "0000101", "0000101", "0001010", "0001001", "0000100", "0000111", "0001000", "0001001", "0001000", "0000101", "0000010", "0000110", "0000010", "0001111", "0001010", "0000110", "0010010", "0010010", "0010001", "0000011", "0001101", "0000110", "0000100", "0001001", "0001011", "0001101", "0001111", "0000110", "0001000", "0000101", "0001010", "0001010", "0000111", "0001000", "0001011", "0000100", "0000011", "0000110", "0001100", "0001010", "0001111", "0001010", "0001001", "0000110", "0000110", "0010001", "0000111", "0010110", "0010010", "0001101", "0001000", "0000101", "0010010", "0010011", "0001100", "0010010", "0010000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000101", "0000101", "0000110", "0000100", "0000100", "0000011", "0001110", "0000011", "0001000", "0000011", "0000101", "0000011", "0001000", "0001011", "0001001", "0000110", "0000100", "0000111", "0001010", "0000111", "0000111", "0000100", "0000001", "0000101", "0000010", "0000010", "0000011", "0001011", "0001100", "0000001", "0000111", "0000010", "0000010", "0000001", "0000010", "0000001", "0000100", "0000110", "0000110", "0010010", "0001111", "0000110", "0001100", "0001101", "0001110", "0001101", "0001001", "0000100", "0001011", "0000011", "0010001", "0001100", "0001000", "0001100", "0001011", "0001010", "0000101", "0000100", "0000010", "0000001", "0000111", "0000010", "0000010", "0000011", "0000001", "0000010", "0000101", "0001010", "0001010", "0000111", "0001000", "0001011", "0000100", "0000110", "0000110", "0001011", "0001011", "0001111", "0001010", "0001010", "0001010", "0000110", "0010001", "0001000", "0001101", "0001100", "0001001", "0001100", "0000010", "0000100", "0000100", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000100", "0000010", "0000111", "0000000", "0000100", "0000010", "0000001", "0000011", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0001100", "0001011", "0000001", "0000111", "0000100", "0000011", "0000011", "0000100", "0000101", "0000010", "0000011", "0000100", "0000110", "0000101", "0000010", "0000100", "0000100", "0000101", "0000101", "0000011", "0000001", "0000011", "0000001", "0000100", "0000011", "0000010", "0000011", "0000011", "0000011", "0000010", "0000011", "0000001", "0000001", "0000111", "0000101", "0000101", "0001100", "0000101", "0000111", "0000001", "0000010", "0000010", "0000001", "0000001", "0000011", "0000001", "0000010", "0000001", "0000010", "0000010", "0000100", "0000001", "0000010", "0000100", "0000001", "0000010", "0000001", "0000110", "0000001", "0000110", "0000100", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000101", "0000011", "0000100", "0001100", "0000111", "0001101", "0000011", "0000010", "0000010", "0000001", "0000001", "0000001", "0000101", "0000010", "0000111", "0000001", "0000011", "0000010", "0000010", "0000011", "0000010", "0000011", "0000001", "0000010", "0000011", "0000010", "0000100", "0000101", "0000001", "0000101", "0001000", "0001000", "0001010", "0010101", "0010011", "0001010", "0010100", "0011000", "0010100", "0001101", "0010000", "0010100", "0000001", "0000001", "0000001", "0000110", "0000101", "0000010", "0000100", "0000100", "0000101", "0000101", "0000011", "0000001", "0000011", "0000001", "0001011", "0000111", "0000100", "0001110", "0001110", "0001101", "0000010", "0001010", "0000101", "0000011", "0001001", "0001010", "0001100", "0010100", "0001000", "0001010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000010", "0000001", "0000001", "0000010", "0000011", "0000001", "0000010", "0000100", "0000001", "0000001", "0000001", "0000110", "0000001", "0000101", "0000100", "0000001", "0000010", "0000011", "0000011", "0000101", "0000100", "0001010", "0000110", "0001000", "0010011", "0001100", "0010110", "0001000", "0001010", "0001010", "0000110", "0000111", "0000110", "0001011", "0000110", "0001011", "0000101", "0000111", "0000101", "0001110", "0001001", "0010000", "0001101", "0001000", "0001110", "0010001", "0001100", "0000110", "0010010", "0000101", "0010011", "0010010", "0010011", "0010101", "0010111", "0010011", "0001101", "0001110", "0001110", "0001100", "0000101", "0000111", "0001000", "0000011", "0000100", "0000100", "0001111", "0001101", "0000101", "0001010", "0001011", "0001100", "0001100", "0000111", "0000011", "0001001", "0000011", "0010001", "0001100", "0000111", "0010000", "0001111", "0001110", "0000101", "0001010", "0000100", "0000011", "0001001", "0001010", "0001011", "0010000", "0000111", "0001010", "0000010", "0000101", "0000101", "0000100", "0000100", "0000110", "0000010", "0000101", "0000011", "0000101", "0000110", "0001001", "0000101", "0000101", "0001001", "0000100", "0001001", "0000100", "0010000", "0001100", "0001011", "0001011", "0000101", "0010000", "0010000", "0001110", "0010100", "0010001", "0001001", "0000100", "0000110", "0001110", "0001000", "0001101", "0000110", "0000110", "0000111", "0000101", "0000101", "0000100", "0001011", "0000101", "0001001", "0000011", "0000111", "0000100", "0001001", "0001000", "0001001", "0001010", "0000101", "0001001", "0001100", "0001000", "0000110", "0000110", "0000010", "0000111", "0000100", "0000100", "0000101", "0001100", "0001100", "0000100", "0001001", "0000111", "0000101", "0000011", "0000110", "0000110", "0000100", "0000101", "0000110", "0001101", "0001011", "0000101", "0001001", "0001001", "0001011", "0001010", "0000111", "0000011", "0000111", "0000010", "0001110", "0001011", "0000110", "0001011", "0001100", "0001011", "0000100", "0000100", "0000010", "0000010", "0000111", "0000010", "0000011", "0000011", "0000001", "0000010", "0000101", "0001100", "0001011", "0001001", "0001001", "0001100", "0000101", "0000100", "0000111", "0001110", "0001100", "0010001", "0001011", "0001011", "0001000", "0000111", "0010011", "0001001", "0010110", "0010100", "0001110", "0001001", "0000101", "0010000", "0010001", "0001011", "0010001", "0001111", "0000100", "0000010", "0000010", "0000011", "0000011", "0000010", "0000100", "0000011", "0000100", "0000010", "0000010", "0000011", "0000011", "0000011", "0000111", "0000010", "0001000", "0000100", "0000100", "0000010", "0000101", "0000111", "0000011", "0000100", "0000101", "0000100", "0000011", "0000110", "0000010", "0000111", "0000110", "0000110", "0001000", "0001111", "0001110", "0000110", "0001001", "0001010", "0001000", "0000011", "0000110", "0000101", "0000100", "0000101", "0000110", "0000100", "0000100", "0000010", "0000011", "0000011", "0000100", "0000100", "0000010", "0000001", "0000011", "0000001", "0000011", "0000101", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000010", "0000011", "0000010", "0000001", "0000100", "0001000", "0001000", "0000110", "0000110", "0001001", "0000100", "0000010", "0000101", "0001010", "0001010", "0001100", "0001000", "0001000", "0000101", "0000110", "0001110", "0000110", "0001111", "0001011", "0001011", "0000011", "0000010", "0000111", "0000110", "0000100", "0000110", "0000101", "0000100", "0000001", "0000010", "0000011", "0000011", "0000100", "0000100", "0000100", "0000100", "0000011", "0000011", "0000011", "0000011", "0000011", "0000111", "0000010", "0000111", "0000100", "0000101", "0000010", "0000110", "0000111", "0000011", "0000110", "0000111", "0000101", "0000011", "0000110", "0000010", "0000110", "0000110", "0000110", "0000111", "0001110", "0001100", "0000100", "0001001", "0000111", "0000110", "0000101", "0000111", "0001000", "0000010", "0000010", "0000010", "0000100", "0000011", "0000010", "0000011", "0000011", "0000011", "0000100", "0000010", "0000001", "0000010", "0000001", "0000110", "0000110", "0000011", "0001000", "0001000", "0000111", "0000001", "0000101", "0000011", "0000010", "0001000", "0000111", "0000111", "0001000", "0000101", "0000110", "0000001", "0000010", "0000010", "0000010", "0000010", "0000011", "0000001", "0000010", "0000001", "0000011", "0000101", "0000110", "0000010", "0000011", "0000100", "0000010", "0000011", "0000010", "0001011", "0000011", "0001000", "0000011", "0000001", "0000010", "0000010", "0000010", "0000011", "0000011", "0001000", "0000101", "0000111", "0010011", "0001011", "0010011", "0000100", "0000101", "0000101", "0000011", "0000100", "0000100", "0000111", "0000011", "0001000", "0000010", "0001001", "0000100", "0000111", "0000101", "0000111", "0000110", "0000100", "0000110", "0000111", "0000101", "0000100", "0000111", "0000010", "0001001", "0000111", "0000110", "0001011", "0001111", "0001101", "0000111", "0001100", "0001101", "0001011", "0000100", "0000110", "0000111", "0000011", "0000100", "0000100", "0001001", "0001000", "0000100", "0000110", "0000111", "0001000", "0000111", "0000100", "0000010", "0000101", "0000010", "0001010", "0000111", "0000100", "0001000", "0001001", "0001000", "0000011", "0000101", "0000011", "0000010", "0000111", "0000101", "0000110", "0001010", "0000100", "0000101", "0000010", "0000100", "0000100", "0000011", "0000011", "0000101", "0000010", "0000011", "0000011", "0000110", "0000101", "0001001", "0000100", "0000100", "0000110", "0000011", "0001000", "0000011", "0001111", "0001001", "0001011", "0000111", "0000011", "0001011", "0001100", "0001010", "0010000", "0001110", "0010001", "0000111", "0001010", "0011111", "0010000", "0011110", "0000101", "0000110", "0000111", "0000100", "0000100", "0000100", "0000110", "0000100", "0001000", "0000011", "0001010", "0000011", "0001000", "0000101", "0001010", "0001000", "0000101", "0001000", "0001011", "0000111", "0000100", "0001010", "0000011", "0001011", "0001001", "0001010", "0001100", "0010011", "0001111", "0001000", "0001011", "0001100", "0001010", "0000110", "0001010", "0001011", "0000011", "0000100", "0000101", "0001000", "0000111", "0000011", "0000101", "0000110", "0000111", "0000110", "0000100", "0000010", "0000101", "0000001", "0001010", "0000110", "0000100", "0001001", "0001000", "0001001", "0000010", "0000110", "0000011", "0000010", "0000111", "0000101", "0000101", "0001001", "0000100", "0000101", "0000111", "0001101", "0001101", "0001010", "0001010", "0001110", "0000110", "0000011", "0001000", "0010001", "0001101", "0010100", "0001110", "0001101", "0000111", "0001001", "0010111", "0001010", "0011110", "0011010", "0010011", "0000110", "0000111", "0010111", "0011000", "0010100", "0011110", "0011001", "0100010", "0010000", "0011001", "0111110", "0100000", "0111111", "0000111", "0001001", "0001001", "0000101", "0000111", "0000110", "0001010", "0000101", "0001010", "0000100", "0001011", "0000100", "0001100", "0000111", "0001110", "0001011", "0000111", "0001011", "0010000", "0001010", "0000101", "0001101", "0000100", "0001110", "0010000", "0001111", "0010001", "0011100", "0010110", "0001111", "0010110", "0011010", "0010110", "0001100", "0001111", "0010100", "0001000", "0001011", "0001011", "0001100", "0001010", "0000101", "0001000", "0001001", "0001010", "0001001", "0000110", "0000011", "0000111", "0000010", "0010001", "0001100", "0000111", "0010100", "0010010", "0010001", "0000011", "0001111", "0000110", "0000101", "0001101", "0010001", "0010011", "0100111", "0010001", "0010110", "0001110", "0011001", "0011100", "0010011", "0010110", "0011101", "0001011", "0000100", "0010001", "0100000", "0011100", "0101010", "0011010", "0011011", "0001101", "0010001", "0101111", "0010100", "0111011", "0110100", "0101001", "0001001", "0010000", "0110100", "0110011", "0101100", "0111101", "0110110", "0001110", "0000111", "0001011", "0010010", "0001010", "0010011", "0010001", "0010100", "0010101", "0001101", "0001110", "0001100", "0101010", "0001100", "0010011", "0001010", "0010010", "0001001", "0011101", "0011101", "0100001", "0011001", "0010001", "0011011", "0100011", "0011001", "0010011", "0100011", "0001010", "0100111", "0100100", "0100110", "0110000", "0110010", "0100111", "0011101", "0100101", "0110010", "0101001", "0010001", "0010110", "0011011", "0010001", "0010110", "0011010", "0110100", "0101110", "0010010", "0100011", "0100111", "0101010", "0100100", "0011011", "0001011", "0011110", "0001001", "1000011", "0101100", "0011100", "1000011", "1000100", "1000000", "0001111", "0101010", "0010100", "0001110", "0011001", "0100111", "0101100", "0111110", "0011010", "0100010", "0001111", "0100000", "0011111", "0011001", "0011001", "0100001", "0001101", "0010000", "0010011", "0101001", "0100000", "0101110", "0100000", "0011111", "0011110", "0010101", "0110100", "0011001", "0110111", "0110001", "0101000", "0100111", "0001011", "0100101", "0101001", "0010110", "0100001", "0011101", "0010011", "0001001", "0001101", "0011010", "0001110", "0011101", "0001111", "0010101", "0010100", "0001101", "0001110", "0001100", "0100111", "0001100", "0010010", "0001011", "0010000", "0001001", "0011100", "0011100", "0011110", "0011000", "0010001", "0011100", "0100101", "0011000", "0010100", "0011010", "0001000", "0011101", "0010100", "0010101", "0011000", "0011001", "0010100", "0001100", "0010010", "0010110", "0010010", "0001101", "0010010", "0010110", "0001010", "0001111", "0001111", "0110000", "0101100", "0010001", "0011101", "0100100", "0101011", "0100110", "0011010", "0001100", "0011100", "0001001", "0110110", "0100100", "0010111", "0101110", "0101110", "0101011", "0001110", "0011100", "0001100", "0001001", "0010101", "0011110", "0100001", "0101101", "0010100", "0011010", "0000110", "0001011", "0001010", "0001000", "0001000", "0001100", "0000101", "0010000", "0000111", "0001110", "0001011", "0010100", "0001011", "0001100", "0011101", "0001000", "0010100", "0001000", "0011011", "0010100", "0010101", "0100010", "0000110", "0010011", "0010100", "0010001", "0011000", "0010110", "0100011", "0010000", "0011001", "1001000", "0100110", "1001000", "0010111", "0011011", "0011110", "0010011", "0010100", "0010001", "1000011", "0010001", "0011001", "0010000", "0010110", "0001100", "0101010", "0110010", "0101101", "0100101", "0011001", "0100111", "0110011", "0100011", "0100011", "0101011", "0001101", "0110000", "0110110", "0110101", "1000011", "1010001", "0111100", "0101110", "0101010", "0110101", "0101101", "0101010", "0110100", "1000001", "0011110", "0100110", "0101101", "1010111", "1001010", "0011111", "0111100", "1000000", "1001001", "1000000", "0101101", "0010100", "0110001", "0001111", "1101011", "1000111", "0101101", "1101000", "1101000", "1100001", "0011010", "0111011", "0011010", "0010100", "0011101", "0101011", "0110010", "1100010", "0101000", "0110110", "0010110", "0110001", "0110000", "0100011", "0100101", "0110010", "0010100", "0011011", "0011110", "0111010", "0110010", "1001000", "0110000", "0101111", "0110000", "0100000", "1010011", "0100100", "1011100", "1010111", "0111101", "0111101", "0010111", "1001110", "1010001", "0111010", "1010000", "1000110", "0001111", "0001000", "0001101", "0011010", "0001110", "0011001", "0101011", "0110101", "0110011", "0100010", "0100111", "0100000", "0100100", "0100000", "0101110", "0011100", "0101001", "0010111", "1001100", "0011011", "1010111", "1000001", "0101101", "1000110", "1011101", "0111110", "0010010", "1010001", "0011000", "1011000", "0111100", "0111101", "1001001", "1001100", "0111010", "0101100", "1000001", "1011011", "1001001", "0010111", "0100000", "0100110", "0001101", "0010001", "0010010", "0101110", "0101000", "0010001", "0011111", "0100100", "0100110", "0100010", "0011010", "0001100", "0011110", "0001001", "0110100", "0100011", "0010110", "0100101", "0100011", "0100011", "0001101", "0010111", "0001010", "0001000", "0001111", "0010011", "0010111", "0011011", "0001110", "0001111", "0001101", "0011001", "0011011", "0010011", "0010011", "0011101", "0001100", "0001110", "0010000", "0100001", "0011010", "0110001", "0011010", "0011001", "0100010", "0010001", "0101111", "0010100", "0111110", "0101010", "0110000", "0100001", "0001001", "0100001", "0100000", "0010110", "0100011", "0011101", "0001111", "0000110", "0001100", "0010000", "0001010", "0010000", "0011010", "0011110", "0100000", "0010110", "0010110", "0010110", "0010111", "0010011", "0011011", "0010001", "0110110", "0001101", "0101011", "0010010", "0110001", "0100101", "0011010", "0101011", "0111000", "0100110", "0001100", "0101111", "0001111", "0110100", "0101001", "0101000", "0110001", "0111001", "0101011", "0100001", "0101101", "1000111", "0110000", "0010100", "0011010", "0100001", "0001011", "0001110", "0010001", "0011110", "0011100", "0001110", "0010101", "0010110", "0011001", "0010111", "0010000", "0001000", "0010011", "0000110", "0100101", "0011010", "0010000", "0100000", "0100000", "0100010", "0001001", "0010011", "0001001", "0000111", "0001110", "0010011", "0011000", "0011101", "0010000", "0010000", "0001000", "0010001", "0010000", "0001101", "0001101", "0010001", "0001001", "0001010", "0001010", "0010100", "0010010", "0101110", "0001110", "0001111", "0100101", "0001010", "0011100", "0001100", "1000010", "0011101", "0111111", "0010110", "0001000", "0010101", "0010111", "0010010", "0011001", "0011000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000101", "0000000", "0000101", "0001010", "0000101", "0000101", "0000000", "0000101", "0000101", "0001010", "0000101", "0000101", "0000000", "0000000", "0000000", "0000000", "0001010", "0000000", "0010100", "0000000", "0001010", "0000000", "0001111", "0000000", "0000000", "0000000", "0000000", "0000101", "0000000", "0000000", "0000000", "0000000", "0000000", "0001010", "0000000", "0000000", "0001010", "0000101", "0001010", "0000101", "0000101", "0000101", "0000000", "0001010", "0001111", "0001010", "0000101", "0010100", "0001010", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000101", "0000101", "0000000", "0001010", "0000101", "0000000", "0000101", "0000000", "0001010", "0001010", "0001111", "0000000", "0000000", "0000101", "0000000", "0000000", "0000101", "0000101", "0000000", "0000101", "0011110", "0001010", "0000101", "0000101", "0000101", "0001010", "0001010", "0000000", "0000000", "0000000", "0010011", "0010101", "0001000", "0010010", "0000111", "0010101", "0001000", "0001011", "0000101", "0010001", "0001101", "0000100", "0011000", "0001101", "0010011", "0001111", "0001000", "0001101", "0010000", "0100101", "0010100", "0001110", "0001101", "0010110", "0001011", "0001101", "0101000", "0000111", "0101001", "0001101", "0010111", "0000110", "0011000", "0010000", "0011000", "0010010", "0010111", "0011101", "0001100", "0001100", "0000110", "0001010", "0001011", "0101100", "0001100", "0001110", "0100001", "0100011", "0110001", "0101000", "0100111", "0101100", "0010110", "0101111", "0011100", "0011011", "0010010", "0101001", "0101000", "0001100", "0001111", "0011011", "0100011", "0101000", "0011000", "0010101", "0010110", "0011010", "0001100", "0010000", "0011101", "0001100", "0010010", "0010111", "0011010", "0001101", "0100111", "0001001", "0100010", "0011000", "0101110", "0001100", "0001001", "0011111", "0010000", "0001011", "0011110", "0100111", "0010110", "0010100", "0101111", "0011010", "0010101", "0011001", "0010100", "0011001", "0010110", "0100011", "0010101", "0100000", "1000011", "1000111", "0011000", "0111111", "0011000", "1000111", "0010001", "0010111", "0001010", "0100111", "0011100", "0001010", "0101000", "0011110", "0101000", "0100011", "0010001", "0011101", "0100010", "0111011", "0101001", "0011110", "0011100", "0110010", "0011001", "0011010", "1000000", "0001111", "0110100", "0010101", "0101110", "0001011", "0101100", "0011010", "0101000", "0011100", "0101100", "0011001", "0010100", "0011011", "0001001", "0010110", "0010001", "1001001", "0010011", "0010110", "0110100", "0111100", "1010000", "0110111", "1000011", "1010000", "0101000", "1000000", "0110110", "0110100", "0100001", "1100001", "1010111", "0011011", "0011001", "0101110", "0111011", "1000110", "1011011", "1001001", "1001111", "1011011", "0101011", "0111011", "0110010", "0010010", "0011101", "0100111", "0101001", "0010011", "0111111", "0001111", "0111000", "0100101", "1001010", "0010101", "0001111", "0110011", "0011001", "0010001", "0100111", "1001000", "0100111", "0100000", "1010100", "0110001", "0101000", "0101000", "0110001", "0111000", "0110010", "0111110", "0100110", "0111010", "0011100", "0011111", "0001011", "0101010", "0010001", "0110000", "0010111", "0100010", "0001110", "0110011", "0100111", "0001110", "0011011", "0101000", "0111001", "0101101", "0011000", "0100101", "0101111", "0101001", "0111000", "0101010", "0100111", "1000101", "0100011", "0100010", "0101010", "0010111", "1000111", "0011110", "1010100", "0010100", "1001100", "0111010", "1011101", "0111001", "1100110", "0110110", "0101111", "1000010", "0010111", "0111000", "0001101", "0110000", "0001101", "0001111", "0100100", "0100111", "0110110", "0100101", "0101101", "0110111", "0011100", "0101110", "0100100", "0100010", "0010100", "0111001", "0110101", "0010000", "0010001", "0100000", "0101000", "0101111", "0100101", "0011110", "0100001", "1000001", "0011101", "0101001", "0100001", "0001100", "0010011", "0011010", "0011100", "0001110", "0101100", "0001010", "0101000", "0011010", "0110011", "0001101", "0001001", "0100011", "0010001", "0001100", "0011010", "0110001", "0011010", "0010101", "0110111", "0100000", "0011010", "0011100", "0011101", "0100001", "0011110", "0101000", "0011000", "0100101", "0101100", "0101110", "0010000", "0100110", "0001111", "0101101", "0011000", "0100001", "0001111", "0110110", "0100110", "0001110", "0010000", "0101001", "0111011", "0101110", "0011000", "0101000", "0110000", "0010111", "0111000", "0101010", "0100110", "1000110", "0100011", "0100001", "0011011", "0010101", "1000000", "0011010", "1000000", "0001111", "0111100", "0100110", "0111010", "0100110", "0111100", "0100001", "0011100", "0100001", "0001100", "0011111", "0001010", "0011100", "0000111", "0001001", "0010100", "0010111", "0011111", "0010110", "0011100", "0011111", "0010000", "0011100", "0011001", "0010111", "0001111", "0101100", "0101001", "0001100", "0001001", "0011100", "0100100", "0101011", "0111010", "0101111", "0110001", "0111001", "0011010", "0100101", "0010101", "0001000", "0001100", "0001111", "0010001", "0001001", "0011000", "0000110", "0010110", "0001110", "0011100", "0001000", "0000110", "0010100", "0001010", "0001010", "0010000", "0011100", "0001111", "0001101", "0100101", "0010110", "0010010", "0010000", "0010111", "0011010", "0010111", "0101000", "0011000", "0100100", "0000101", "0000110", "0000010", "0000101", "0000010", "0000110", "0001000", "0001011", "0000110", "0010001", "0001101", "0000100", "0000001", "0001110", "0010010", "0010000", "0001000", "0001100", "0001111", "0000010", "0010100", "0001100", "0001101", "0010101", "0001100", "0001011", "0000010", "0001001", "0100010", "0001101", "0100110", "0001010", "0100110", "0100000", "0110011", "0100100", "1000011", "0100100", "0011110", "0110100", "0010010", "0101101", "0000111", "0000010", "0000001", "0000010", "0000001", "0000010", "0000110", "0000100", "0000100", "0000010", "0000001", "0001100", "0000010", "0000011", "0000010", "0000101", "0001101", "0000100", "0000001", "0000011", "0000100", "0000100", "0000111", "0000101", "0000110", "0000111", "0000100", "0000101", "0000101", "0000010", "0000001", "0000001", "0000010", "0000011", "0000011", "0000001", "0000010", "0000011", "0000011", "0000001", "0000001", "0000010", "0000001", "0000111", "0000100", "0000010", "0000010", "0000011", "0000100", "0000010", "0000010", "0000001", "0000011", "0000011", "0000011", "0000100", "0000011", "0000111", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000111", "0000001", "0000010", "0000001", "0000001", "0000011", "0000001", "0000000", "0001001", "0000010", "0000010", "0000010", "0000010", "0000001", "0000010", "0001011", "0000100", "0000011", "0000010", "0000011", "0000001", "0000010", "0000111", "0000001", "0000001", "0000010", "0000001", "0000001", "0000100", "0000011", "0000010", "0000001", "0000001", "0001100", "0000001", "0000010", "0000010", "0000010", "0001011", "0000101", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000001", "0000011", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000000", "0000001", "0000000", "0000111", "0000010", "0000001", "0000001", "0000010", "0000011", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000111", "0000001", "0000010", "0000001", "0000000", "0000010", "0000001", "0000000", "0000110", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0001100", "0000011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000001", "0000010", "0000001", "0000001", "0000011", "0000010", "0000010", "0000001", "0000001", "0001100", "0000001", "0000011", "0000010", "0000010", "0001011", "0000100", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000011", "0000010", "0000000", "0000000", "0000001", "0000000", "0000111", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000010", "0000001", "0000000", "0000010", "0000001", "0000000", "0000100", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0001100", "0000011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000111", "0000001", "0000010", "0000010", "0000010", "0001011", "0000101", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000011", "0000000", "0000000", "0000001", "0000000", "0000110", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000010", "0000010", "0000001", "0000010", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000011", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0001011", "0000010", "0000010", "0000001", "0000001", "0000001", "0000000", "0000111", "0000001", "0000010", "0000010", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000110", "0000001", "0000010", "0000011", "0000010", "0001011", "0000100", "0000001", "0000001", "0000010", "0000010", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000011", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000011", "0000000", "0000000", "0000001", "0000000", "0000111", "0000001", "0000000", "0000010", "0000001", "0000010", "0000000", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000011", "0000001", "0000001", "0000001", "0000010", "0000001", "0000000", "0000000", "0000011", "0000010", "0000001", "0000010", "0000000", "0000000", "0000010", "0000001", "0000011", "0000010", "0000000", "0000001", "0000000", "0000111", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000011", "0000010", "0000000", "0000010", "0000001", "0000000", "0000000", "0001011", "0000011", "0000001", "0000001", "0000000", "0000000", "0000000", "0000111", "0000000", "0000010", "0000010", "0000000", "0000000", "0000011", "0000010", "0000010", "0000000", "0000001", "0000100", "0000001", "0000010", "0000100", "0000010", "0001011", "0000111", "0000001", "0000001", "0000011", "0000011", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000011", "0000001", "0000001", "0000001", "0000011", "0000010", "0000001", "0000010", "0000001", "0000001", "0000100", "0000000", "0000000", "0000001", "0000000", "0000111", "0000001", "0000000", "0000011", "0000001", "0000010", "0000000", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000011", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000100", "0000010", "0000010", "0000010", "0000001", "0000001", "0000011", "0000010", "0000100", "0000010", "0000001", "0000010", "0000010", "0000111", "0000010", "0000011", "0000010", "0000001", "0000010", "0000010", "0000000", "0000011", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0001100", "0000011", "0000001", "0000001", "0000001", "0000000", "0000000", "0000111", "0000010", "0000011", "0000011", "0000001", "0000001", "0000011", "0000010", "0000010", "0000010", "0000001", "0000101", "0000001", "0000100", "0000101", "0000010", "0001011", "0000100", "0000001", "0000001", "0000011", "0000011", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000100", "0000001", "0000001", "0000001", "0000100", "0000010", "0000010", "0000010", "0000010", "0000001", "0000110", "0000001", "0000000", "0000010", "0000001", "0000111", "0000001", "0000010", "0000011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000100", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000101", "0000111", "0000100", "0001010", "0001000", "0000011", "0001001", "0001000", "0001011", "0001010", "0000101", "0001000", "0001001", "0001101", "0001101", "0001000", "0000111", "0001101", "0000110", "0000110", "0001111", "0000100", "0001011", "0000101", "0001000", "0000011", "0001000", "0000011", "0000101", "0001101", "0000100", "0000010", "0000001", "0000001", "0000001", "0000001", "0001000", "0010000", "0000101", "0000101", "0001100", "0001100", "0010001", "0001011", "0001110", "0010001", "0001001", "0001101", "0001000", "0001001", "0000111", "0001001", "0001101", "0000100", "0000101", "0000011", "0000101", "0000101", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0001011", "0000100", "0000111", "0001001", "0001010", "0000101", "0001110", "0000100", "0001101", "0001000", "0010000", "0000100", "0000011", "0001011", "0000101", "0000111", "0001000", "0010000", "0001001", "0000111", "0001100", "0000111", "0000110", "0001001", "0000101", "0000101", "0000101", "0000100", "0000010", "0000101", "0001110", "0001111", "0000101", "0001101", "0000101", "0001101", "0000011", "0000100", "0000011", "0000110", "0000101", "0000010", "0001010", "0000101", "0000111", "0000110", "0000011", "0000100", "0000110", "0001111", "0001010", "0000101", "0000101", "0001000", "0000100", "0000100", "0010000", "0000011", "0001010", "0000100", "0001101", "0000011", "0001100", "0001010", "0010000", "0001111", "0010001", "0001001", "0001000", "0001010", "0000011", "0001000", "0000111", "0010001", "0000101", "0000110", "0001110", "0001110", "0010011", "0001101", "0010000", "0010010", "0001001", "0001111", "0001110", "0001110", "0001001", "0010111", "0011001", "0000111", "0000110", "0001101", "0010000", "0010011", "0010010", "0010000", "0010000", "0010001", "0001001", "0001100", "0001100", "0000100", "0000111", "0001001", "0001010", "0000101", "0010000", "0000100", "0001110", "0001001", "0010001", "0000101", "0000011", "0001100", "0000110", "0001000", "0001001", "0010000", "0001001", "0000111", "0010110", "0001101", "0001010", "0001010", "0001100", "0001101", "0001100", "0010000", "0001010", "0001111", "0001111", "0010000", "0000110", "0010010", "0000111", "0010100", "0000100", "0000110", "0000011", "0001001", "0000111", "0000010", "0000100", "0000111", "0001010", "0001000", "0000100", "0000111", "0001000", "0000110", "0001011", "0000111", "0000110", "0001100", "0000110", "0000101", "0000111", "0000011", "0001011", "0000101", "0001001", "0000010", "0001000", "0000101", "0001000", "0001100", "0001001", "0000101", "0000100", "0000111", "0000011", "0000111", "0000111", "0000111", "0000011", "0000011", "0000101", "0000110", "0001000", "0000101", "0000111", "0001000", "0000100", "0000111", "0001000", "0001000", "0000110", "0010001", "0010100", "0000101", "0000011", "0001011", "0001111", "0010000", "0010110", "0010001", "0010010", "0011101", "0001101", "0010001", "0000101", "0000010", "0000011", "0000100", "0000101", "0000011", "0000110", "0000010", "0000101", "0000100", "0001001", "0000010", "0000001", "0000101", "0000010", "0001000", "0000100", "0000111", "0000100", "0000011", "0001101", "0000111", "0000110", "0000100", "0001001", "0001001", "0001001", "0001111", "0001001", "0001110", "0001000", "0001001", "0000011", "0001011", "0000101", "0001101", "0000001", "0000010", "0000011", "0000011", "0000011", "0000001", "0000001", "0000011", "0000011", "0000011", "0000001", "0000010", "0000011", "0000001", "0001000", "0000010", "0000010", "0000100", "0000010", "0000010", "0000001", "0000010", "0000110", "0000010", "0001010", "0000010", "0001001", "0001000", "0001100", "0001111", "0001110", "0000111", "0000110", "0001000", "0000011", "0000111", "0000111", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000010", "0000011", "0000100", "0001100", "0000011", "0000001", "0000101", "0000101", "0000111", "0001100", "0001001", "0001010", "0010001", "0001000", "0001011", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000000", "0000000", "0000001", "0000000", "0000111", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000011", "0000010", "0000010", "0000101", "0000100", "0000101", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000010", "0000011", "0000011", "0000001", "0000001", "0000011", "0000011", "0000011", "0000001", "0000010", "0000011", "0000001", "0001000", "0000010", "0000010", "0000100", "0000010", "0000010", "0000001", "0000001", "0000011", "0000001", "0000010", "0000001", "0000010", "0000010", "0000011", "0001100", "0000110", "0000011", "0000011", "0000110", "0000010", "0000101", "0000111", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000010", "0000010", "0000001", "0001011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000010", "0000001", "0000000", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000000", "0000000", "0000001", "0000000", "0000111", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000011", "0000010", "0000010", "0000001", "0000010", "0000010", "0000010", "0000111", "0000010", "0000010", "0000011", "0000001", "0000010", "0000010", "0000001", "0000100", "0000010", "0000101", "0000001", "0000100", "0000011", "0000100", "0001100", "0000011", "0000010", "0000001", "0000010", "0000001", "0000001", "0000111", "0000010", "0000001", "0000010", "0000010", "0000010", "0000011", "0000010", "0000010", "0000010", "0000001", "0000011", "0000001", "0000010", "0000001", "0000001", "0001011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000011", "0000001", "0000000", "0000010", "0000001", "0000111", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000011", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000010", "0000000", "0000010", "0000010", "0000011", "0000101", "0000101", "0000011", "0000010", "0000011", "0000001", "0000011", "0000011", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000011", "0000110", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000011", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000011", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000010", "0000011", "0000010", "0000010", "0000100", "0000010", "0000010", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000010", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000010", "0000000", "0000001", "0000001", "0000010", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000010", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000000", "0000000", "0000001", "0000000", "0000000", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000010", "0000010", "0000001", "0000010", "0000001", "0000011", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000010", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000001", "0000010", "0000010", "0000011", "0000010", "0000011", "0000100", "0000010", "0000010", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000001", "0000000", "0000000", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000000", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000100", "0000000", "0000001", "0000001", "0000000", "0000001", "0000010", "0000000", "0000010", "0000001", "0000011", "0000001", "0000010", "0000011", "0000100", "0000111", "0000101", "0000011", "0000010", "0000011", "0000001", "0000011", "0000100", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000010", "0000010", "0000010", "0000001", "0000011", "0000111", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000000", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000100", "0000001", "0000010", "0000001", "0000001", "0000011", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000010", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000011", "0000010", "0000001", "0000001", "0000011", "0000011", "0000010", "0000001", "0000010", "0000011", "0000001", "0000111", "0000010", "0000010", "0000100", "0000010", "0000010", "0000010", "0000001", "0000100", "0000010", "0000100", "0000001", "0000100", "0000010", "0000011", "0001100", "0000011", "0000001", "0000001", "0000010", "0000001", "0000001", "0000111", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0001011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000111", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000011", "0000001", "0000011", "0000001", "0000010", "0000010", "0000010", "0000010", "0000001", "0000001", "0000011", "0000011", "0000011", "0000001", "0000010", "0000011", "0000001", "0000111", "0000010", "0000010", "0000011", "0000010", "0000010", "0000001", "0000001", "0000011", "0000001", "0000011", "0000001", "0000010", "0000011", "0000100", "0001100", "0001001", "0000100", "0000100", "0001000", "0000011", "0000110", "0000111", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000010", "0000010", "0000001", "0001011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000100", "0000010", "0000011", "0000001", "0000000", "0000001", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000000", "0000000", "0000001", "0000000", "0000111", "0000001", "0000001", "0000001", "0000001", "0000001", "0000000", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0001010", "0001011", "0000100", "0001101", "0000101", "0001111", "0000010", "0000011", "0000011", "0000100", "0000011", "0000001", "0000001", "0000100", "0000100", "0000011", "0000010", "0000011", "0000100", "0000001", "0001000", "0000011", "0000011", "0000101", "0000011", "0000011", "0000001", "0000011", "0001000", "0000011", "0001011", "0000011", "0001011", "0001000", "0001101", "0001111", "0001100", "0000111", "0000110", "0000111", "0000010", "0000110", "0000111", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000011", "0000010", "0000010", "0000011", "0000110", "0001101", "0000011", "0000001", "0000110", "0000111", "0001001", "0001110", "0001011", "0001100", "0010101", "0001001", "0001100", "0000010", "0000000", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000011", "0000000", "0000000", "0000001", "0000000", "0000111", "0000001", "0000001", "0000001", "0000001", "0000011", "0000010", "0000001", "0000001", "0000100", "0000011", "0000011", "0001000", "0000101", "0000111", "0010001", "0010000", "0000110", "0010011", "0000111", "0010100", "0000100", "0000110", "0000011", "0001000", "0000111", "0000010", "0000110", "0000111", "0001010", "0001000", "0000100", "0000110", "0001000", "0001000", "0001011", "0000111", "0000110", "0001011", "0000110", "0000101", "0001001", "0000011", "0001010", "0000100", "0001000", "0000010", "0000111", "0000101", "0001000", "0001100", "0001011", "0000101", "0000101", "0001001", "0000011", "0001000", "0000111", "0001010", "0000011", "0000100", "0000111", "0001000", "0001011", "0000111", "0001010", "0001010", "0000101", "0001000", "0001001", "0001001", "0000110", "0010100", "0010101", "0000110", "0000011", "0001101", "0001111", "0010011", "0010111", "0010011", "0010010", "0011100", "0001110", "0010010", "0000111", "0000010", "0000100", "0000101", "0000110", "0000011", "0001000", "0000010", "0000111", "0000101", "0001010", "0000011", "0000010", "0000111", "0000011", "0001000", "0000101", "0001001", "0000101", "0000100", "0001111", "0001000", "0000111", "0000101", "0001010", "0001011", "0001010", "0001111", "0001010", "0001111", "0001011", "0001100", "0000100", "0001000", "0000100", "0001010", "0000011", "0000101", "0000011", "0000111", "0000101", "0000010", "0001011", "0000110", "0000111", "0000110", "0000011", "0000101", "0000110", "0010000", "0001011", "0000101", "0000101", "0001001", "0000101", "0000100", "0010001", "0000100", "0001011", "0000101", "0001110", "0000100", "0001101", "0001010", "0001111", "0001111", "0001111", "0001000", "0000111", "0001000", "0000011", "0000110", "0001000", "0010010", "0000101", "0000110", "0001110", "0001111", "0010100", "0001101", "0010010", "0010101", "0001010", "0001111", "0001110", "0001110", "0001001", "0011000", "0011000", "0000111", "0000111", "0001011", "0001111", "0010000", "0001111", "0001100", "0001110", "0001110", "0000110", "0001001", "0001101", "0000101", "0000111", "0001010", "0001011", "0000101", "0010001", "0000100", "0001110", "0001001", "0010011", "0000101", "0000100", "0001101", "0000110", "0001000", "0001010", "0010010", "0001010", "0001000", "0010110", "0001101", "0001010", "0001010", "0001100", "0001101", "0001100", "0001111", "0001000", "0001110", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000100", "0000110", "0000100", "0001001", "0000111", "0000011", "0000111", "0000111", "0001010", "0001001", "0000100", "0000111", "0001000", "0001011", "0001100", "0000111", "0000111", "0001100", "0000110", "0000101", "0001100", "0000011", "0001001", "0000100", "0000101", "0000010", "0000101", "0000010", "0000011", "0001100", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0001000", "0001100", "0000100", "0000101", "0001001", "0001010", "0001101", "0001001", "0001011", "0001101", "0000111", "0001011", "0000110", "0000111", "0000110", "0000101", "0001101", "0000100", "0000100", "0000010", "0000011", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0001001", "0000011", "0000110", "0000111", "0001000", "0000100", "0001011", "0000011", "0001011", "0000110", "0001101", "0000100", "0000011", "0001000", "0000101", "0000111", "0000111", "0001100", "0000111", "0000101", "0001001", "0000101", "0000100", "0000111", "0000100", "0000011", "0000011", "0000010", "0000010", "0000100", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000011", "0000010", "0000001", "0000010", "0000000", "0000001", "0000010", "0000001", "0000011", "0000010", "0000001", "0000010", "0000001", "0000111", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000000", "0000011", "0000001", "0000001", "0000010", "0000001", "0000000", "0000001", "0001100", "0000011", "0000001", "0000001", "0000001", "0000000", "0000000", "0000111", "0000001", "0000011", "0000010", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000001", "0000101", "0000001", "0000011", "0000101", "0000010", "0001100", "0000100", "0000001", "0000001", "0000011", "0000011", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000100", "0000001", "0000001", "0000001", "0000011", "0000010", "0000001", "0000010", "0000001", "0000001", "0000101", "0000000", "0000000", "0000001", "0000000", "0000111", "0000001", "0000001", "0000011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000010", "0000010", "0000001", "0000010", "0000000", "0000000", "0000010", "0000001", "0000011", "0000010", "0000000", "0000001", "0000000", "0000111", "0000001", "0000001", "0000000", "0000000", "0000001", "0000001", "0000000", "0000011", "0000010", "0000000", "0000010", "0000001", "0000000", "0000000", "0001011", "0000011", "0000001", "0000001", "0000000", "0000000", "0000000", "0000111", "0000000", "0000010", "0000010", "0000000", "0000000", "0000011", "0000010", "0000010", "0000000", "0000001", "0000100", "0000001", "0000010", "0000100", "0000010", "0001011", "0000111", "0000001", "0000001", "0000010", "0000011", "0000000", "0000000", "0000001", "0000001", "0000000", "0000000", "0000011", "0000001", "0000001", "0000001", "0000011", "0000010", "0000001", "0000010", "0000001", "0000001", "0000100", "0000000", "0000000", "0000001", "0000000", "0000111", "0000010", "0000000", "0000011", "0000001", "0000010", "0000000", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000011", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000010", "0000010", "0000001", "0000010", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000010", "0000001", "0000000", "0000001", "0000001", "0000000", "0000011", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0001011", "0000011", "0000010", "0000001", "0000001", "0000001", "0000000", "0000111", "0000001", "0000010", "0000010", "0000000", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000110", "0000001", "0000010", "0000011", "0000010", "0001011", "0000100", "0000001", "0000001", "0000010", "0000010", "0000001", "0000000", "0000001", "0000001", "0000000", "0000000", "0000011", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000001", "0000011", "0000000", "0000000", "0000001", "0000000", "0000111", "0000001", "0000000", "0000010", "0000010", "0000010", "0000000", "0000001", "0000001", "0000010", "0000001", "0000001", "0000000", "0000001", "0000011", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000010", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000010", "0000001", "0000000", "0000010", "0000001", "0000000", "0000100", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0001100", "0000011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000001", "0000010", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0001000", "0000001", "0000011", "0000010", "0000010", "0001100", "0000101", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000011", "0000000", "0000000", "0000001", "0000000", "0000110", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000000", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000111", "0000001", "0000010", "0000001", "0000000", "0000011", "0000001", "0000000", "0000111", "0000010", "0000001", "0000010", "0000010", "0000001", "0000001", "0001011", "0000011", "0000010", "0000001", "0000001", "0000001", "0000001", "0000111", "0000001", "0000001", "0000010", "0000001", "0000001", "0000011", "0000010", "0000010", "0000001", "0000001", "0001100", "0000001", "0000010", "0000010", "0000010", "0001011", "0000101", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000001", "0000010", "0000010", "0000010", "0000001", "0000001", "0000011", "0000010", "0000000", "0000000", "0000001", "0000000", "0000111", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000001", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000100", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000010", "0000001", "0000011", "0000000", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000010", "0000001", "0000110", "0000001", "0000010", "0000001", "0000001", "0000011", "0000001", "0000001", "0001001", "0000011", "0000010", "0000010", "0000011", "0000010", "0000011", "0001100", "0000111", "0000101", "0000011", "0000110", "0000010", "0000101", "0000110", "0000001", "0000001", "0000010", "0000000", "0000001", "0000101", "0000011", "0000011", "0000001", "0000001", "0001011", "0000001", "0000010", "0000010", "0000010", "0001100", "0000100", "0000001", "0000010", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000001", "0000011", "0000001", "0000001", "0000001", "0000001", "0000011", "0000010", "0000001", "0000001", "0000010", "0000010", "0000001", "0000000", "0000001", "0000000", "0000111", "0000010", "0000001", "0000001", "0000010", "0000011", "0000001", "0000001", "0000001", "0000010", "0000001", "0000010", "0000001", "0000001", "0000101", "0001010", "0001010", "0000011", "0001010", "0000100", "0001101", "0001101", "0010010", "0001000", "0011101", "0010101", "0001000", "0000010", "0010111", "0011111", "0011010", "0001101", "0010110", "0011010", "0000011", "0011111", "0010111", "0010110", "0100111", "0010011", "0010011", "0000100", "0001111", "0110001", "0010011", "0111010", "0001110", "0110110", "0101101", "1000111", "0101101", "1011000", "0101101", "0100111", "0111010", "0010101", "0110100", "0000111", "0000100", "0000001", "0000011", "0000010", "0000011", "0000111", "0000101", "0000101", "0000100", "0000010", "0001101", "0000011", "0000100", "0000011", "0001000", "0001101", "0000101", "0000010", "0000110", "0000111", "0001000", "0001100", "0001010", "0001010", "0010001", "0001000", "0001011", "0000101", "0000010", "0000010", "0000010", "0000011", "0000011", "0000100", "0000001", "0000011", "0000011", "0000100", "0000010", "0000001", "0000011", "0000001", "0000111", "0000100", "0000011", "0000011", "0000011", "0000111", "0000011", "0000011", "0000010", "0000100", "0000101", "0000101", "0000111", "0000101", "0001001", "0101101", "0110001", "0010000", "0101111", "0010010", "0110110", "0010100", "0011100", "0001101", "0101110", "0100001", "0001100", "0010101", "0100010", "0110011", "0101000", "0010101", "0100001", "0101001", "0100000", "0110010", "0100011", "0100000", "0111010", "0011111", "0011011", "0100011", "0010001", "0110110", "0010110", "0110100", "0001100", "0110001", "0011111", "0101111", "0100000", "0110000", "0011101", "0010111", "0100101", "0001101", "0011111", "0001011", "0100110", "0001010", "0001100", "0011100", "0011110", "0101010", "0011110", "0100100", "0101010", "0010110", "0100100", "0100001", "0011110", "0010100", "0111010", "0110110", "0010000", "0001101", "0100001", "0101011", "0110010", "0111011", "0110000", "0110100", "1000111", "0100001", "0101101", "0011011", "0001010", "0010000", "0010101", "0010110", "0001100", "0100011", "0001000", "0011111", "0010100", "0100111", "0001011", "0001000", "0011011", "0001110", "0001011", "0010101", "0100110", "0010101", "0010000", "0110001", "0011101", "0010111", "0010101", "0011110", "0100001", "0011110", "0101101", "0011011", "0101001", "0100001", "0100010", "0001100", "0100111", "0010000", "0101111", "0011011", "0100111", "0010000", "0111100", "0101101", "0010001", "0011010", "0101110", "1000001", "0110100", "0011100", "0101011", "0110110", "0100101", "1000000", "0110000", "0101101", "1001111", "0101000", "0100111", "0101000", "0011011", "1010011", "0100010", "1011010", "0010110", "1010101", "0111110", "1100010", "0111110", "1100111", "0110110", "0110000", "1000010", "0010111", "0111001", "0001100", "0101101", "0001101", "0001101", "0100000", "0100110", "0110010", "0100010", "0101010", "0110011", "0011001", "0101101", "0100010", "0100000", "0010011", "0110110", "0110000", "0010000", "0010000", "0011111", "0100111", "0101110", "0110000", "0100110", "0101000", "0111011", "0011011", "0100110", "0100000", "0001100", "0010001", "0011000", "0011011", "0001101", "0101000", "0001001", "0100011", "0011000", "0110000", "0001101", "0001001", "0100000", "0010000", "0001100", "0011000", "0101100", "0010111", "0010100", "0110100", "0011110", "0011001", "0011010", "0011001", "0011111", "0011011", "0101010", "0011001", "0100110", "0111110", "1000010", "0010110", "0110101", "0010100", "0111010", "0001101", "0010010", "0001000", "0011100", "0010101", "0001000", "0101011", "0010110", "0011111", "0011011", "0001101", "0010110", "0011010", "0111111", "0011111", "0010111", "0010101", "0100110", "0010100", "0010100", "1000101", "0001011", "0101010", "0010001", "0100011", "0001001", "0100001", "0010011", "0011101", "0010110", "0100110", "0010110", "0010001", "0010000", "0000101", "0001011", "0010010", "1001111", "0010101", "0010111", "0111000", "0111111", "1010101", "0111011", "1001001", "1010110", "0101011", "1000100", "0111010", "0111000", "0100100", "1011000", "1010000", "0011001", "0011010", "0110100", "1000010", "1001110", "1010000", "1000010", "1000110", "1001100", "0100100", "0110001", "0110100", "0010010", "0100000", "0101010", "0101100", "0010101", "1000011", "0010001", "0111100", "0101001", "1001111", "0010110", "0010000", "0110111", "0011100", "0010010", "0101001", "1001100", "0101001", "0100010", "1011011", "0110101", "0101100", "0101011", "0101101", "0110100", "0101111", "1000100", "0101010", "0111110");
  constant classconst : class_sim := (1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4);
  
  SIGNAL start_bit_int	                       	  	  		: STD_LOGIC; 
  --Random Value Generation Signals
  SIGNAL clock_val							: STD_LOGIC_VECTOR(127 DOWNTO 0);
  SIGNAL seed_ready                       	  		  	: STD_LOGIC;  
  SIGNAL out_ready_int                               			: STD_LOGIC;
  SIGNAL out_val_int                      	  		  	: STD_LOGIC;  
  SIGNAL out_int							: STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL out_buffer							: STD_LOGIC_VECTOR(2879 DOWNTO 0);
  
  --Position and Level Hypervector Generation Signals
  SIGNAL index							        : integer range 0 to 2880;
  SIGNAL full_HV							: integer range 0 to 91;
  SIGNAL pos_HV_num							: integer range 0 to 76;
  --SIGNAL	pos_HVs							: vector_of_std_logic_vector2880(0 TO 74)  := (others => (others => '0')); 
  SIGNAL	posHV_data						: STD_LOGIC_VECTOR(2879 DOWNTO 0);
  SIGNAL	posHV_out						: STD_LOGIC_VECTOR(2879 DOWNTO 0);
  SIGNAL posHV_Wen		                    	  		: STD_LOGIC;
  SIGNAL posHV_Ren		                    	  		: STD_LOGIC;
  SIGNAL posHV_slv					           	: STD_LOGIC_VECTOR(6 DOWNTO 0);
  SIGNAL lev_HV_num							: integer range 0 to 117;
  SIGNAL lev_buffer							: STD_LOGIC_VECTOR(2879 DOWNTO 0); 
  --SIGNAL	lev_HVs							: vector_of_std_logic_vector2880(0 TO 116)  := (others => (others => '0'));   
  SIGNAL	levHV_data						: STD_LOGIC_VECTOR(2879 DOWNTO 0);
  SIGNAL	levHV_out						: STD_LOGIC_VECTOR(2879 DOWNTO 0);
  SIGNAL levHV_Wen		                    	  		: STD_LOGIC;
  SIGNAL levHV_Ren		                    	  		: STD_LOGIC;
  SIGNAL levHV_slv					           	: STD_LOGIC_VECTOR(6 DOWNTO 0);
 
  --Memory signals
  SIGNAL bins_addr_in             					: STD_LOGIC_VECTOR (14 DOWNTO 0) := "000000000000000";
  SIGNAL bins_rom_out                 					: STD_LOGIC_VECTOR (6 DOWNTO 0) := "0000000";
  
  --Division signals
  --SIGNAL divisor						        : STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000001010000";
  --SIGNAL dividend						        : STD_LOGIC_VECTOR(31 DOWNTO 0);
  --SIGNAL divres					           	: STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
  --SIGNAL div_flag		                    	  		: std_logic_vector(0 downto 0) := "0"; 


  
  --Class training counter
  SIGNAL class_HV_num							: integer range 0 to 5; 
  --Class testing counter
  SIGNAL test_HV_num							: integer range 0 to 5; 


  --Sample Encode counters
  SIGNAL enc_bin_num							: STD_LOGIC_VECTOR (6 DOWNTO 0) := "0000000";
  SIGNAL enc_sample_num							: integer range 0 to 80;  
  --Encode Values
  SIGNAL bin_value							: integer range 0 to 116;
  SIGNAL pos_val							: STD_LOGIC_VECTOR(2879 DOWNTO 0);
  SIGNAL lev_val							: STD_LOGIC_VECTOR(2879 DOWNTO 0);
  SIGNAL res_vec							: STD_LOGIC_VECTOR(2879 DOWNTO 0);
  --SIGNAL res_total							: STD_LOGIC_VECTOR(31 DOWNTO 0);
  

  
  --Retrain signals
  --SIGNAL retrain_diff							: STD_LOGIC_VECTOR(31 DOWNTO 0);
  --SIGNAL retrain_int_val						: STD_LOGIC_VECTOR(31 DOWNTO 0);
  --SIGNAL diff_slv						        : STD_LOGIC_VECTOR(31 DOWNTO 0);
  --SIGNAL divres_retrain			           	     	: STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
  
  --Result Signals
  SIGNAL done_bit_int	                    	  		  	: STD_LOGIC;
  SIGNAL correct_cnt_slv						: STD_LOGIC_VECTOR(6 DOWNTO 0); 
  SIGNAL total_cnt_slv							: STD_LOGIC_VECTOR(6 DOWNTO 0);
  SIGNAL hexone								: STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL hextwo								: STD_LOGIC_VECTOR (6 DOWNTO 0);
  
 

BEGIN

--Memory, Division instantiations
	--Bins
  ROMinst:    		Bins_ROM					PORT MAP(bins_addr_in,CLOCK_50,bins_rom_out);
	--RNG
  Xoshinst: 		rng_xoshiro128plusplus 				PORT MAP(CLOCK_50,RESET,seed_ready,clock_val,out_ready_int,out_val_int,out_int);
  
	--Div for classes
  --Divinst: 			lpmDiv							PORT MAP(CLOCK_50,divisor,dividend,divres);
  
	--Div for retrain
  --retrainOne: 		lpmDiv							PORT MAP(CLOCK_50,divisor,diff_slv,divres_retrain);

	--Storing level and pos HVs
  posHVs_inst:    posHV_RAM						PORT MAP(CLOCK_50,posHV_data,posHV_slv,posHV_Ren,posHV_slv,posHV_Wen,posHV_out);
  levHVs_inst:    levHV_RAM						PORT MAP(CLOCK_50,levHV_data,levHV_slv,levHV_Ren,levHV_slv,levHV_Wen,levHV_out);
		
--HDC Process		
  HDC_Aud: Process(CLOCK_50,RESET)
  
  
  
  variable classOne								: class_vector := (others => (others => '0'));   
  variable classTwo								: class_vector := (others => (others => '0'));   
  variable classThree								: class_vector := (others => (others => '0'));   
  variable classFour								: class_vector := (others => (others => '0'));  
  variable classOneTrained							: class_vector := (others => (others => '0'));   
  variable classTwoTrained							: class_vector := (others => (others => '0'));   
  variable classThreeTrained							: class_vector := (others => (others => '0'));   
  variable classFourTrained							: class_vector := (others => (others => '0'));  
  variable testMX								: class_vector := (others => (others => '0'));  
 
    --Class vectors
  --variable class_one_total							: STD_LOGIC_VECTOR(31 DOWNTO 0);
  --variable class_two_total							: STD_LOGIC_VECTOR(31 DOWNTO 0);
  --variable class_three_total							: STD_LOGIC_VECTOR(31 DOWNTO 0);
  --variable class_four_total							: STD_LOGIC_VECTOR(31 DOWNTO 0);
  
    --Inference vars
  variable diff_one								: STD_LOGIC_VECTOR(31 DOWNTO 0);
  variable diff_two								: STD_LOGIC_VECTOR(31 DOWNTO 0);
  variable diff_three								: STD_LOGIC_VECTOR(31 DOWNTO 0);
  variable diff_four								: STD_LOGIC_VECTOR(31 DOWNTO 0);
  
  
  variable prediction								: integer range 1 to 4; 
  variable sample_class								: integer range 1 to 4; 
  variable res_total								: STD_LOGIC_VECTOR(31 DOWNTO 0);
  variable testnum								: integer range 0 to 80;
  
  
  
  BEGIN

  				--Reset 
				if (RESET = '1') then
					clock_val 				<= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
					start_bit_int				<= '0';
					seed_ready				<= '0';
					out_ready_int 				<= '0';
					out_buffer				<= (others => '0');

					index					<= 0;
					full_HV					<= 0;
					pos_HV_num				<= 0;
					--pos_HVs				<= (others => (others => '0')); 
					posHV_data				<= (others => '0');
					posHV_Wen	 			<= '0';
					posHV_Ren	 			<= '0';
					posHV_slv				<= "0000000";
					lev_HV_num				<= 0;
					lev_buffer				<= (others => '0');
					--lev_HVs				<= (others => (others => '0')); 
					levHV_data				<= (others => '0');
					levHV_Wen	 			<= '0';
					levHV_Ren	 			<= '0';
					levHV_slv				<= "0000000";
					
					bins_addr_in				<= "000000000000000";

					--divisor				<= "00000000000000000000000001010000";
					--dividend				<= "00000000000000000000000000000000";
					--div_flag				<= "0";

					class_HV_num				<= 0;
					--class_one_total			:= "00000000000000000000000000000000";
					--class_two_total			:= "00000000000000000000000000000000";
					--class_three_total			:= "00000000000000000000000000000000";
					--class_four_total			:= "00000000000000000000000000000000";

					enc_bin_num				<= "0000000";
					enc_sample_num				<= 0;
					bin_value 				<= 0;
					pos_val					<= (others => '0');
					lev_val					<= (others => '0');
					res_vec					<= (others => '0');
					res_total				:= "00000000000000000000000000000000";

					test_HV_num				<= 0;
					diff_one				:= "00000000000000000000000000000000";
					diff_two				:= "00000000000000000000000000000000";
					diff_three				:= "00000000000000000000000000000000";
					diff_four				:= "00000000000000000000000000000000";
					
					--retrain_diff				<= "00000000000000000000000000000000";
					--retrain_int_val			<= "00000000000000000000000000000000";
					--diff_slv				<= "00000000000000000000000000000000";
					
					done_bit_int				<= '0';
					correct_cnt_slv 			<= "0000000";
					total_cnt_slv 				<= "0000000";
					
					testnum					:= 0;
					prediction 				:= 1;
					sample_class				:= 1;
					hexone					<= "1111111";
					hextwo					<= "1111111";
					
					classOne				:= (others => (others => '0')); 
					classTwo				:= (others => (others => '0')); 
					classThree				:= (others => (others => '0')); 
					classFour				:= (others => (others => '0')); 
					classOneTrained				:= (others => (others => '0')); 
					classTwoTrained				:= (others => (others => '0')); 
					classThreeTrained			:= (others => (others => '0')); 
					classFourTrained			:= (others => (others => '0')); 
					testMX					:= (others => (others => '0')); 
					
					Mealy_state 		<= START;
			
  
  
  			elsif(RISING_EDGE(CLOCK_50)) then  
				clock_val 		<= clock_val + "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
				IF (clock_val  = "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111") then  
					clock_val 	<= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
				end if;

	  --User flips switch to start HDC process
	  			CASE Mealy_State IS
				WHEN START =>
					IF SW = '1' then  			
						start_bit_int <= '1';
						Mealy_state <= POSITION_HVS;
					ELSE
						Mealy_state <= START;  		-- wait until user ready and presses button
					END IF;
					  
		--Position HVs generation
				WHEN POSITION_HVS =>
					IF(pos_HV_num < 75) then
						Mealy_state 				<= HV_SETUP;
					ELSE
						posHV_Wen				<= '0';
						Mealy_state 				<= LEV_HV_FIRST;
					END IF;

					
				WHEN HV_SETUP =>
					IF(full_HV < 90) then
						IF (out_val_int = '1') then
							out_ready_int 		<= '1';
							index 				<= to_integer(to_unsigned(full_HV,128) * 32);					
							Mealy_state			<= HV_STORE;
						ELSE
							Mealy_state			<= HV_SETUP;
						END IF;
					ELSE
						Mealy_state 		<= HV_READY;
					END IF;
					
					
				WHEN HV_STORE =>	
				 	out_buffer((index + 31) DOWNTO (index)) <= out_int;
					full_HV 						<= full_HV + 1;
					Mealy_state 						<= HV_SETUP;
					
				WHEN HV_READY =>
					IF (pos_HV_num = 74) then
							--pos_HVs(pos_HV_num)	<= out_buffer;
							posHV_Wen				<= '1';
							posHV_data				<= out_buffer;
							posHV_slv				<= posHV_slv + "0000001";
							full_HV 				<= 0;
							pos_HV_num 				<= pos_HV_num + 1;
							Mealy_state 				<= POSITION_HVS;
					ELSE
							--pos_HVs(pos_HV_num)	<= out_buffer;
							posHV_Wen				<= '1';
							posHV_data				<= out_buffer;
							posHV_slv				<= posHV_slv + "0000001";
							full_HV 				<= 0;
							pos_HV_num 				<= pos_HV_num + 1;
							Mealy_state 				<= POSITION_HVS;
					END IF;
					
					
				WHEN LEV_HV_FIRST =>
					IF(lev_HV_num < 1) then
						IF(full_HV < 90) then
							IF (out_val_int = '1') then
								out_ready_int 				<= '1';
								index 					<= to_integer(to_unsigned(full_HV,128) * 32);
								out_buffer((index + 31) DOWNTO (index)) <= out_int;
								full_HV 				<= full_HV + 1;
							END IF;
						ELSIF (full_HV = 90) then
							--lev_HVs(0)				<= out_buffer;
							levHV_Wen				<= '1';
							levHV_data				<= out_buffer;
							levHV_slv				<= levHV_slv + "0000001";
							lev_HV_num 				<= 1;
							full_HV 				<= 0;
						END IF;
					ELSE
						index 		<= 0;
						Mealy_state 	<= LEVEL_HVS;
					END IF;
					
				WHEN LEVEL_HVS =>
					IF(lev_HV_num < 117) then
						--lev_buffer 				<= lev_HVs(lev_HV_num - 1);
						lev_buffer 				<= levHV_data;
						index 					<= to_integer(to_unsigned(lev_HV_num - 1,128) * 24);
						Mealy_state 				<= LEVEL_HV_FLIP; 
					ELSE
						levHV_Wen				<= '0';
						Mealy_state 				<= AUDIO_ENC; 
					END IF;
					
				WHEN LEVEL_HV_FLIP =>
						
						lev_buffer((index + 23) DOWNTO (index)) <= not lev_buffer((index + 23) DOWNTO (index));
						Mealy_state 			<= LEVEL_HV_SET; 
					
				WHEN LEVEL_HV_SET =>
						levHV_Wen				<= '1';
						levHV_data				<= lev_buffer;
						levHV_slv				<= levHV_slv + "0000001";
						lev_HV_num 				<= lev_HV_num + 1;
						Mealy_state 				<= LEVEL_HVS;
				
				WHEN AUDIO_ENC =>
					levHV_Ren						<= '1';
					posHV_Ren						<= '1';
					IF (class_HV_num = 4) then
						Mealy_state 				<= AUDIO_ENC_TEST;
					ELSIF (enc_sample_num < 80) then
						
						IF (enc_bin_num = "1001011") then
							enc_sample_num 			<= enc_sample_num + 1; --increasing sample number so reset bins addr to sample
							
							IF (class_HV_num = 0) then
								bins_addr_in 				<= std_logic_vector(to_unsigned(enc_sample_num,15)); 
							ELSIF (class_HV_num = 1) then
								bins_addr_in 				<= std_logic_vector(to_unsigned(enc_sample_num,15)) + "001110101001100"; 
							ELSIF (class_HV_num = 2) then
								bins_addr_in 				<= std_logic_vector(to_unsigned(enc_sample_num,15)) + "011101010011000"; 
							ELSE 
								bins_addr_in 				<= std_logic_vector(to_unsigned(enc_sample_num,15)) + "101011111100100"; 
							END IF;
							
							enc_bin_num 				<= "0000000";
							Mealy_state 				<= AUDIO_ENC;
						ELSE
							Mealy_state 				<= ENC_BIN_SETUP; 
						END IF;
					ELSE
						Mealy_state 				<= TRAIN; 
					END IF;
				
				WHEN ENC_BIN_SETUP =>
						posHV_slv 					<= enc_bin_num;
						---------------------------------------
						--real impl
						levHV_slv 					<= bins_rom_out;
						--sim impl
						--levHV_slv					<= binsconst(to_integer(unsigned(bins_addr_in)));
						---------------------------------------
						Mealy_state 				<= ENC_BIN_SET; 
				
				WHEN ENC_BIN_SET =>
						pos_val					<= posHV_out;
						lev_val					<= levHV_out;
						Mealy_state 				<= ENC_BIN_VAL; 
						
				WHEN ENC_BIN_VAL =>
						res_vec					<= pos_val AND lev_val;
						enc_bin_num 				<= enc_bin_num + "0000001"; --increasing bin so need to add 100 to addr
						bins_addr_in				<= bins_addr_in + "000000001100100";						
						Mealy_state 				<= TRAIN; 
				
				
				--this becomes the new train
				WHEN TRAIN =>
					--this or separate state
				IF(class_HV_num < 4) then
					for I in 2879 downto 0 loop
						IF (res_vec(I) = '1') then
							IF(class_HV_num = 0) then
								classOne(I) := classOne(I) + "0000001";
									IF(classOne(I) = "1010000") then --if reaches 80, add one to trained 
										classOneTrained(I) := classOneTrained(I) + "0000001";
										classOne(I) :=  "0000000";
									ELSE
									END IF;
							ELSIF(class_HV_num = 1) then
								classTwo(I) := classTwo(I) + "0000001";
									IF(classTwo(I) = "1010000") then --if reaches 80, add one to trained 
										classTwoTrained(I) := classTwoTrained(I) + "0000001";
										classTwo(I) :=  "0000000";
									ELSE
									END IF;
							ELSIF(class_HV_num = 2) then
								classThree(I) := classThree(I) + "0000001";
									IF(classThree(I) = "1010000") then --if reaches 80, add one to trained 
										classThreeTrained(I) := classThreeTrained(I) + "0000001";
										classThree(I) :=  "0000000";
									ELSE
									END IF;
							ELSE
								classFour(I) := classFour(I) + "0000001";
									IF(classFour(I) = "1010000") then --if reaches 80, add one to trained
										classFourTrained(I) := classFourTrained(I) + "0000001";
										classFour(I) :=  "0000000";
									ELSE
									END IF;
							END IF;
							--res_total				:= res_total + "00000000000000000000000000000001";
						ELSE
						END IF;
					end loop;	
					IF (enc_sample_num = 80) THEN
						enc_sample_num <= 0;
						class_HV_num <= class_HV_num + 1;
					ELSE
					END IF;
					Mealy_state 				<= AUDIO_ENC; 
				ELSE
				Mealy_state 				<= AUDIO_ENC_TEST; 
				END IF;

	
				WHEN AUDIO_ENC_TEST =>	
					IF(test_HV_num < 4) THEN
						IF(enc_sample_num < 20) THEN
							IF (enc_bin_num = "1001011") then
								IF (test_HV_num = 0) then
									bins_addr_in 				<= std_logic_vector(to_unsigned(enc_sample_num,15)) + "000000001010000"; --+80
								ELSIF (test_HV_num = 1) then
									bins_addr_in 				<= std_logic_vector(to_unsigned(enc_sample_num,15)) + "001110110011100"; --7500+80
								ELSIF (test_HV_num = 2) then
									bins_addr_in 				<= std_logic_vector(to_unsigned(enc_sample_num,15)) + "011101011101000"; --15000+80
								ELSE
									bins_addr_in 				<= std_logic_vector(to_unsigned(enc_sample_num,15)) + "101100000110100"; --22500+80
								END IF;
								Mealy_state 				<= INF;
							ELSE
								posHV_slv 					<= enc_bin_num;
								--------------------------------------
								--real impl
								levHV_slv 					<= bins_rom_out;
								--sim impl
								--levHV_slv					<= binsconst(to_integer(unsigned(bins_addr_in)));
								---------------------------------------
								--might not need the read enables
								levHV_Ren						<= '1';
								posHV_Ren						<= '1';
								
								IF(levHV_Ren = '1' AND posHV_Ren = '1') then
									pos_val						<= posHV_out;
									lev_val						<= levHV_out;
								ELSE
									Mealy_state 					<= AUDIO_ENC;
								END IF;
								
								res_vec						<= pos_val AND lev_val;
								
								MEALY_STATE					<= TEST_BIN_VEC;

							END IF;
						ELSE
							enc_sample_num <= 0;
							test_HV_num 	<= test_HV_num + 1;
						END IF;
					ELSE
						Mealy_state 				<= RESULT;
					END IF;

			WHEN TEST_BIN_VEC =>
											--this or separate state
				for I in 2879 downto 0 loop
					IF (res_vec(I) = '1') then
						testMX(I) := testMX(I) + "0000001";
					ELSE
					END IF;
				end loop;	
				
				enc_bin_num 				<= enc_bin_num + "0000001";
				bins_addr_in				<= bins_addr_in + "000000001100100";
				Mealy_state 				<= AUDIO_ENC_TEST; 
				
		
				WHEN INF =>
					enc_bin_num 				<= "0000000";
					------------------------------------------
					--for sim
					sample_class				:= classconst(testnum);
					testnum 						:= testnum + 1;
					------------------------------------------
					for J in 3 downto 0 loop
						-- have to check which is greater for each index because no abs
							for I in 2879 downto 0 loop
								IF (J = 0) then
									IF (testMX(I) > classOneTrained(I)) then
										diff_one := testMX(I) - classOneTrained(I) + diff_one;
									ELSE
										diff_one := classOneTrained(I) - testMX(I) + diff_one;
									END IF;
								ELSIF (J = 1) then
									IF (testMX(I) > classTwoTrained(I)) then
										diff_two := testMX(I) - classTwoTrained(I) + diff_two;
									ELSE
										diff_two := classTwoTrained(I) - testMX(I) + diff_two;
									END IF;
								ELSIF (J = 2) then
									IF (testMX(I) > classThreeTrained(I)) then
										diff_three := testMX(I) - classThreeTrained(I) + diff_three;
									ELSE
										diff_three := classThreeTrained(I) - testMX(I) + diff_three;
									END IF;
								ELSE	
									IF (testMX(I) > classFourTrained(I)) then
										diff_four := testMX(I) - classFourTrained(I) + diff_four;
									ELSE
										diff_four := classFourTrained(I) - testMX(I) + diff_four;
									END IF;
								END IF;
							end loop;	
					end loop;
					
					IF((diff_one < diff_two	) AND (diff_one < diff_three) AND (diff_one < diff_four)) then
						prediction 					:= 1;
--						retrain_diff				<= diff_one;
					ELSIF((diff_two	 < diff_three) AND (diff_two	 < diff_four)) then
						prediction 					:= 2;
--						retrain_diff				<= diff_two;
					ELSIF((diff_three < diff_four)) then
						prediction 					:= 3;
--						retrain_diff				<= diff_three;
					ELSE 
						prediction 					:= 4;
--						retrain_diff				<= diff_four;
					END IF;
--						--diff_slv						<= std_logic_vector(to_unsigned(retrain_diff,32));
--						diff_slv						<= retrain_diff;
						total_cnt_slv 				<= total_cnt_slv + "0000001";
						enc_sample_num				<= enc_sample_num + 1;
						Mealy_state 				<= INF_RES;
					--need to know sample class to know if need to retrain
					
					
					
				WHEN INF_RES =>
					testMX					:= (others => (others => '0')); 
					diff_one				:= "00000000000000000000000000000000";
					diff_two				:= "00000000000000000000000000000000";
					diff_three				:= "00000000000000000000000000000000";
					diff_four				:= "00000000000000000000000000000000";
					IF (prediction = sample_class) then
						Mealy_state 				<= AUDIO_ENC_TEST;
						correct_cnt_slv 			<= correct_cnt_slv + "0000001";
						--res_total					:= "00000000000000000000000000000000";
					ELSE
						Mealy_state 				<= RETRAIN;
						--res_total					:= "00000000000000000000000000000000";
					END IF;
					

--check for overflow
				WHEN RETRAIN =>
					for I in 2879 downto 0 loop
						IF(prediction = 1) THEN
							IF(classOneTrained(I) > 1) THEN
								classOneTrained(I)			:= classOneTrained(I) - "0000001";
							ELSE
							END IF;
						ELSIF(prediction = 2) THEN
							IF(classTwoTrained(I) > 1) THEN
								classTwoTrained(I)			:= classTwoTrained(I) - "0000001";
							ELSE
							END IF;
						ELSIF(prediction = 3) THEN
							IF(classThreeTrained(I) > 1) THEN
								classThreeTrained(I)			:= classThreeTrained(I) - "0000001";
							ELSE
							END IF;
						ELSE
							IF(classFourTrained(I) > 1) THEN
								classFourTrained(I)			:= classFourTrained(I) - "0000001";
							ELSE
							END IF;
						END IF;	
						
						
						IF(sample_class = 1) then
							IF(classOneTrained(I) < 126) THEN
								classOneTrained(I)			:= classOneTrained(I) + "0000001";
							ELSE
							END IF;
						ELSIF(sample_class = 2) then
							IF(classTwoTrained(I) < 126) THEN
								classTwoTrained(I)			:= classTwoTrained(I) + "0000001";
							ELSE
							END IF;
						ELSIF(sample_class = 3) then
							IF(classThreeTrained(I) < 126) THEN
								classThreeTrained(I)			:= classThreeTrained(I) + "0000001";
							ELSE
							END IF;
						ELSE 
							IF(classFourTrained(I) < 126) THEN
								classFourTrained(I)			:= classFourTrained(I) + "0000001";
							ELSE
							END IF;
						END IF;
					end loop;
--from retain, loop back to Audio enc and do the next sample
					Mealy_state 				<= AUDIO_ENC_TEST;

					

				
				WHEN RESULT =>
					IF(correct_cnt_slv = "0000000") then  --0
						hexone					<= "1111111";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0000001") then --1
						hexone					<= "1001111";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0000010") then --2
						hexone					<= "0010010";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0000011") then --3
						hexone					<= "0000110";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0000100") then --4
						hexone					<= "1001100";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0000101") then --5
						hexone					<= "0100100";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0000110") then --6
						hexone					<= "0100000";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0000111") then --7
						hexone					<= "0001111";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0001000") then --8
						hexone					<= "0000000";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0001001") then --9
						hexone					<= "0001100";
						hextwo					<= "1111111";
					ELSIF(correct_cnt_slv = "0001010") then --10
						hexone					<= "0000001";
						hextwo					<= "0110000";
					ELSIF(correct_cnt_slv = "0001011") then --11
						hexone					<= "1001111";
						hextwo					<= "1001111";
					ELSIF(correct_cnt_slv = "0001100") then --12
						hexone					<= "0010010";
						hextwo					<= "1001111";
					ELSIF(correct_cnt_slv = "0001101") then --13
						hexone					<= "0000110";
						hextwo					<= "1001111";
					ELSIF(correct_cnt_slv = "0001110") then --14
						hexone					<= "1001100";
						hextwo					<= "1001111";
					ELSIF(correct_cnt_slv = "0001111") then --15
						hexone					<= "0100100";
						hextwo					<= "1001111";
					ELSIF(correct_cnt_slv = "0010000") then --16
						hexone					<= "0100000";
						hextwo					<= "1001111";
					ELSIF(correct_cnt_slv = "0010001") then --17
						hexone					<= "0001111";
						hextwo					<= "1001111";
					ELSIF(correct_cnt_slv = "0010010") then --18
						hexone					<= "0000000";
						hextwo					<= "1001111";
					ELSIF(correct_cnt_slv = "0010011") then --19
						hexone					<= "0001100";
						hextwo					<= "1001111";
					ELSIF(correct_cnt_slv = "0010100") then --20
						hexone					<= "0000001";
						hextwo					<= "0010010";
					ELSIF(correct_cnt_slv = "0010101") then --21
						hexone					<= "1001111";
						hextwo					<= "0010010";
					ELSIF(correct_cnt_slv = "0010110") then --22
						hexone					<= "0010010";
						hextwo					<= "0010010";
					ELSIF(correct_cnt_slv = "0010101") then --23
						hexone					<= "0000110";
						hextwo					<= "0010010";
					ELSIF(correct_cnt_slv = "0010110") then --24
						hexone					<= "1001100";
						hextwo					<= "0010010";
					ELSIF(correct_cnt_slv = "0010111") then --25
						hexone					<= "0100100";
						hextwo					<= "0010010";
					ELSIF(correct_cnt_slv = "0011000") then --26
						hexone					<= "0100000";
						hextwo					<= "0010010";	
					ELSIF(correct_cnt_slv = "0011001") then --27
						hexone					<= "0001111";
						hextwo					<= "0010010";		
					ELSIF(correct_cnt_slv = "0011010") then --28
						hexone					<= "0000000";
						hextwo					<= "0010010";
					ELSIF(correct_cnt_slv = "0011011") then --29
						hexone					<= "0001100";
						hextwo					<= "0010010";
					ELSIF(correct_cnt_slv = "0011100") then --30
						hexone					<= "0000001";
						hextwo					<= "0000110";						
					ELSIF(correct_cnt_slv = "0011101") then --31
						hexone					<= "1001111";
						hextwo					<= "0000110";		
					ELSIF(correct_cnt_slv = "0011110") then --32
						hexone					<= "0010010";
						hextwo					<= "0000110";	
					ELSIF(correct_cnt_slv = "0011111") then --33
						hexone					<= "0000110";
						hextwo					<= "0000110";	
					ELSIF(correct_cnt_slv = "0100000") then --34
						hexone					<= "1001100";
						hextwo					<= "0000110";
					ELSIF(correct_cnt_slv = "0100001") then --35
						hexone					<= "0100100";
						hextwo					<= "0000110";
					ELSIF(correct_cnt_slv = "0100010") then --36
						hexone					<= "0100000";
						hextwo					<= "0000110";						
					ELSIF(correct_cnt_slv = "0100011") then --37
						hexone					<= "0001111";
						hextwo					<= "0000110";	
					ELSIF(correct_cnt_slv = "0100100") then --38
						hexone					<= "0000000";
						hextwo					<= "0000110";							
					ELSIF(correct_cnt_slv = "0100101") then --39
						hexone					<= "0001100";
						hextwo					<= "0000110";							
					ELSIF(correct_cnt_slv = "0100110") then --40
						hexone					<= "0000001";
						hextwo					<= "1001100";		
					ELSIF(correct_cnt_slv = "0100111") then --41
						hexone					<= "1001111";
						hextwo					<= "1001100";								
					ELSIF(correct_cnt_slv = "0101000") then --42
						hexone					<= "0010010";
						hextwo					<= "1001100";								
					ELSIF(correct_cnt_slv = "0101001") then --43
						hexone					<= "0000110";
						hextwo					<= "1001100";							
					ELSIF(correct_cnt_slv = "0101010") then --44
						hexone					<= "1001100";
						hextwo					<= "1001100";	
					ELSIF(correct_cnt_slv = "0101011") then --45
						hexone					<= "0100100";
						hextwo					<= "1001100";	
					ELSIF(correct_cnt_slv = "0101100") then --46
						hexone					<= "0100000";
						hextwo					<= "1001100";	
					ELSIF(correct_cnt_slv = "0101101") then --47
						hexone					<= "0001111";
						hextwo					<= "1001100";	
					ELSIF(correct_cnt_slv = "0101110") then --48
						hexone					<= "0000000";
						hextwo					<= "1001100";	
					ELSIF(correct_cnt_slv = "0101111") then --49
						hexone					<= "0001100";
						hextwo					<= "1001100";
					ELSIF(correct_cnt_slv = "0110000") then --50
						hexone					<= "0000001";
						hextwo					<= "0100100";
					ELSIF(correct_cnt_slv = "0110001") then --51
						hexone					<= "1001111";
						hextwo					<= "0100100";
					ELSIF(correct_cnt_slv = "0110010") then --52
						hexone					<= "0010010";
						hextwo					<= "0100100";
					ELSIF(correct_cnt_slv = "0110011") then --53
						hexone					<= "0000110";
						hextwo					<= "0100100";
					ELSIF(correct_cnt_slv = "0110100") then --54
						hexone					<= "1001100";
						hextwo					<= "0100100";
					ELSIF(correct_cnt_slv = "0110101") then --55
						hexone					<= "0100100";
						hextwo					<= "0100100";
					ELSIF(correct_cnt_slv = "0110110") then --56
						hexone					<= "0100000";
						hextwo					<= "0100100";
					ELSIF(correct_cnt_slv = "0110111") then --57
						hexone					<= "0001111";
						hextwo					<= "0100100";						
					ELSIF(correct_cnt_slv = "0111000") then --58
						hexone					<= "0000000";
						hextwo					<= "0100100";	
					ELSIF(correct_cnt_slv = "0111001") then --59
						hexone					<= "0001100";
						hextwo					<= "0100100";	
					ELSIF(correct_cnt_slv = "0111010") then --60
						hexone					<= "0000001";
						hextwo					<= "0100000";	
					ELSIF(correct_cnt_slv = "0111011") then --61
						hexone					<= "1001111";
						hextwo					<= "0100000";	
					ELSIF(correct_cnt_slv = "0111100") then --62
						hexone					<= "0010010";
						hextwo					<= "0100000";
					ELSIF(correct_cnt_slv = "0111101") then --63
						hexone					<= "0000110";
						hextwo					<= "0100000";
					ELSIF(correct_cnt_slv = "0111110") then --64
						hexone					<= "1001100";
						hextwo					<= "0100000";						
					ELSIF(correct_cnt_slv = "0111111") then --65
						hexone					<= "0100100";
						hextwo					<= "0100000";		
					ELSIF(correct_cnt_slv = "1000000") then --66
						hexone					<= "0100000";
						hextwo					<= "0100000";	
					ELSIF(correct_cnt_slv = "1000001") then --67
						hexone					<= "0001111";
						hextwo					<= "0100000";	
					ELSIF(correct_cnt_slv = "1000010") then --68
						hexone					<= "0000000";
						hextwo					<= "0100000";						
					ELSIF(correct_cnt_slv = "1000011") then --69
						hexone					<= "0001100";
						hextwo					<= "0100000";								
					ELSIF(correct_cnt_slv = "1000100") then --70
						hexone					<= "0000001";
						hextwo					<= "0001111";							
					ELSIF(correct_cnt_slv = "1000101") then --71
						hexone					<= "1001111";
						hextwo					<= "0001111";
					ELSIF(correct_cnt_slv = "1000110") then --72
						hexone					<= "0010010";
						hextwo					<= "0001111";
					ELSIF(correct_cnt_slv = "1000111") then --73
						hexone					<= "0000110";
						hextwo					<= "0001111";
					ELSIF(correct_cnt_slv = "1001000") then --74
						hexone					<= "1001100";
						hextwo					<= "0001111";
					ELSIF(correct_cnt_slv = "1001001") then --75
						hexone					<= "0100100";
						hextwo					<= "0001111";						
					ELSIF(correct_cnt_slv = "1001010") then --76
						hexone					<= "0100000";
						hextwo					<= "0001111";								
					ELSIF(correct_cnt_slv = "1001011") then --77
						hexone					<= "0001111";
						hextwo					<= "0001111";		
					ELSIF(correct_cnt_slv = "1001100") then --78
						hexone					<= "0000000";
						hextwo					<= "0001111";							
					ELSIF(correct_cnt_slv = "1001101") then --79
						hexone					<= "0001100";
						hextwo					<= "0001111";	
					ELSE
						hexone					<= "0000001";
						hextwo					<= "0000000";	
					END IF;
					done_bit_int				<= '1';
					Mealy_state 				<= RESULT;
				END CASE;	
				
			end if;
  END PROCESS HDC_Aud;
	 START_BIT  <= start_bit_int;
	 DONE_BIT	<= done_bit_int;
	 CORRECT_HEXONE <= hexone;
	 CORRECT_HEXTWO <= hextwo;
--  PRED_LIGHT <= PRED_LIGHT_INT;
--  DONE_LIGHT <= IDLE_LIGHT;
END Behavior;
